* SPICE3 file created from mult_32.ext - technology: sky130A

X0 net101 clknet_1_0__leaf__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND clknet_1_0__leaf__0461_ net101 VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 net101 clknet_1_0__leaf__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR clknet_1_0__leaf__0461_ net101 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 net61 _0985_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 _0985_/a_891_413# _0985_/a_193_47# _0985_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X6 _0985_/a_561_413# _0985_/a_27_47# _0985_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7 VPWR net71 _0985_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 net61 _0985_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X9 _0985_/a_381_47# _0083_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VGND _0985_/a_634_159# _0985_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X11 VPWR _0985_/a_891_413# _0985_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X12 _0985_/a_466_413# _0985_/a_193_47# _0985_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X13 VPWR _0985_/a_634_159# _0985_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.17887 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X14 _0985_/a_634_159# _0985_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X15 _0985_/a_634_159# _0985_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.17887 ps=1.26 w=0.75 l=0.15
X16 _0985_/a_975_413# _0985_/a_193_47# _0985_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VGND _0985_/a_1059_315# _0985_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X18 _0985_/a_193_47# _0985_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 _0985_/a_891_413# _0985_/a_27_47# _0985_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X20 _0985_/a_592_47# _0985_/a_193_47# _0985_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X21 VPWR _0985_/a_1059_315# _0985_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X22 _0985_/a_1017_47# _0985_/a_27_47# _0985_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X23 _0985_/a_193_47# _0985_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 _0985_/a_466_413# _0985_/a_27_47# _0985_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X25 VGND _0985_/a_891_413# _0985_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X26 _0985_/a_381_47# _0083_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 VGND net71 _0985_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X28 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=707.2962 ps=6.62772k w=0.87 l=1.05
X29 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=450.85931 ps=4.80461k w=0.55 l=1.05
X30 VPWR _0243_ _0770_/a_382_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X31 _0770_/a_297_47# control0.add _0770_/a_79_21# VGND sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X32 _0770_/a_297_47# _0243_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 VGND _0389_ _0770_/a_297_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X34 VPWR _0770_/a_79_21# _0390_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X35 _0770_/a_79_21# control0.add VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X36 _0770_/a_382_297# _0389_ _0770_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X37 VGND _0770_/a_79_21# _0390_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X38 net82 clknet_1_0__leaf__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X39 VGND clknet_1_0__leaf__0459_ net82 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X40 net82 clknet_1_0__leaf__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X41 VPWR clknet_1_0__leaf__0459_ net82 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X42 VPWR net34 _0968_/a_193_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X43 _0968_/a_193_297# control0.state\[1\] _0968_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X44 _0486_ control0.state\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X45 VGND net34 _0486_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X46 _0968_/a_109_297# control0.state\[0\] _0486_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X47 VGND control0.state\[0\] _0486_ VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X48 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X49 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X50 VPWR acc0.A\[6\] _0822_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X51 VGND acc0.A\[6\] _0430_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X52 _0822_/a_109_297# net64 _0430_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X53 _0430_ net64 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X54 _0753_/a_465_47# _0233_ _0753_/a_381_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X55 VGND _0375_ _0753_/a_561_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X56 VPWR _0231_ _0753_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X57 _0753_/a_297_297# _0233_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X58 _0753_/a_297_297# _0375_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X59 VPWR _0222_ _0753_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X60 _0753_/a_381_47# _0222_ _0753_/a_79_21# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.18362 ps=1.215 w=0.65 l=0.15
X61 _0753_/a_297_297# _0343_ _0753_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X62 VPWR _0753_/a_79_21# _0377_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X63 _0753_/a_79_21# _0343_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.18362 pd=1.215 as=0.16087 ps=1.145 w=0.65 l=0.15
X64 VGND _0753_/a_79_21# _0377_ VGND sky130_fd_pr__nfet_01v8 ad=0.16087 pd=1.145 as=0.169 ps=1.82 w=0.65 l=0.15
X65 _0753_/a_561_47# _0231_ _0753_/a_465_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X66 VPWR net55 _0684_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X67 _0316_ _0684_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X68 VGND net55 _0684_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X69 _0684_/a_59_75# acc0.A\[27\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X70 _0316_ _0684_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X71 _0684_/a_145_75# acc0.A\[27\] _0684_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X72 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X73 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X74 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.97
X75 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.97
X76 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X77 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X78 acc0.A\[21\] _1021_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X79 _1021_/a_891_413# _1021_/a_193_47# _1021_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X80 _1021_/a_561_413# _1021_/a_27_47# _1021_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X81 VPWR net107 _1021_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X82 acc0.A\[21\] _1021_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X83 _1021_/a_381_47# _0119_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X84 VGND _1021_/a_634_159# _1021_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X85 VPWR _1021_/a_891_413# _1021_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X86 _1021_/a_466_413# _1021_/a_193_47# _1021_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X87 VPWR _1021_/a_634_159# _1021_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X88 _1021_/a_634_159# _1021_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X89 _1021_/a_634_159# _1021_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X90 _1021_/a_975_413# _1021_/a_193_47# _1021_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X91 VGND _1021_/a_1059_315# _1021_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X92 _1021_/a_193_47# _1021_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X93 _1021_/a_891_413# _1021_/a_27_47# _1021_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X94 _1021_/a_592_47# _1021_/a_193_47# _1021_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X95 VPWR _1021_/a_1059_315# _1021_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X96 _1021_/a_1017_47# _1021_/a_27_47# _1021_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X97 _1021_/a_193_47# _1021_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X98 _1021_/a_466_413# _1021_/a_27_47# _1021_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X99 VGND _1021_/a_891_413# _1021_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X100 _1021_/a_381_47# _0119_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X101 VGND net107 _1021_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X102 VPWR _0281_ _0805_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X103 VPWR _0402_ _0805_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14222 pd=1.335 as=0.06615 ps=0.735 w=0.42 l=0.15
X104 _0805_/a_181_47# _0286_ _0805_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X105 VGND _0402_ _0805_/a_181_47# VGND sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X106 _0805_/a_27_47# _0286_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06615 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X107 _0417_ _0805_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14222 ps=1.335 w=1 l=0.15
X108 _0417_ _0805_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X109 _0805_/a_109_47# _0281_ _0805_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X110 _0736_/a_56_297# _0219_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X111 VPWR _0362_ _0736_/a_56_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X112 _0107_ _0181_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X113 _0736_/a_139_47# _0362_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.2665 ps=2.12 w=0.65 l=0.15
X114 _0736_/a_311_297# _0363_ _0736_/a_56_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X115 _0107_ _0181_ _0736_/a_311_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X116 VGND _0363_ _0107_ VGND sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X117 _0107_ _0219_ _0736_/a_139_47# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X118 VPWR _0226_ _0598_/a_382_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.305 ps=2.61 w=1 l=0.15
X119 _0598_/a_297_47# _0229_ _0598_/a_79_21# VGND sky130_fd_pr__nfet_01v8 ad=0.3705 pd=3.74 as=0.169 ps=1.82 w=0.65 l=0.15
X120 _0598_/a_297_47# _0226_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X121 VGND _0227_ _0598_/a_297_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X122 VPWR _0598_/a_79_21# _0230_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.28 ps=2.56 w=1 l=0.15
X123 _0598_/a_79_21# _0229_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.15
X124 _0598_/a_382_297# _0227_ _0598_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X125 VGND _0598_/a_79_21# _0230_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X126 VPWR acc0.A\[13\] _0299_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X127 _0299_ acc0.A\[13\] _0667_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X128 _0667_/a_113_47# net40 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X129 _0299_ net40 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X130 VPWR clknet_0__0459_ clkbuf_1_0__f__0459_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X131 VPWR clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X132 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X133 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X134 VPWR clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X135 VPWR clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X136 clkbuf_1_0__f__0459_/a_110_47# clknet_0__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X137 clkbuf_1_0__f__0459_/a_110_47# clknet_0__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X138 VGND clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X139 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X140 VGND clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X141 clkbuf_1_0__f__0459_/a_110_47# clknet_0__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X142 VGND clknet_0__0459_ clkbuf_1_0__f__0459_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X143 VGND clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X144 VPWR clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X145 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X146 VGND clknet_0__0459_ clkbuf_1_0__f__0459_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X147 VGND clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X148 VPWR clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X149 VGND clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X150 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X151 clkbuf_1_0__f__0459_/a_110_47# clknet_0__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X152 VPWR clknet_0__0459_ clkbuf_1_0__f__0459_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X153 VPWR clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X154 VPWR clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X155 VGND clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X156 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X157 VGND clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X158 VGND clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X159 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X160 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X161 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X162 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X163 VPWR clkbuf_1_0__f__0459_/a_110_47# clknet_1_0__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X164 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X165 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X166 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X167 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X168 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X169 clknet_1_0__leaf__0459_ clkbuf_1_0__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
X170 VPWR _0121_ hold30/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X171 VGND hold30/a_285_47# hold30/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.5
X172 net177 hold30/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X173 VGND _0121_ hold30/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X174 VPWR hold30/a_285_47# hold30/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.5
X175 hold30/a_285_47# hold30/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X176 hold30/a_285_47# hold30/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X177 net177 hold30/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X178 VPWR acc0.A\[10\] hold41/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X179 VGND hold41/a_285_47# hold41/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X180 net188 hold41/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X181 VGND acc0.A\[10\] hold41/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X182 VPWR hold41/a_285_47# hold41/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X183 hold41/a_285_47# hold41/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X184 hold41/a_285_47# hold41/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X185 net188 hold41/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X186 VPWR acc0.A\[24\] hold52/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X187 VGND hold52/a_285_47# hold52/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X188 net199 hold52/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X189 VGND acc0.A\[24\] hold52/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X190 VPWR hold52/a_285_47# hold52/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X191 hold52/a_285_47# hold52/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X192 hold52/a_285_47# hold52/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X193 net199 hold52/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X194 VPWR acc0.A\[25\] hold63/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X195 VGND hold63/a_285_47# hold63/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X196 net210 hold63/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X197 VGND acc0.A\[25\] hold63/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X198 VPWR hold63/a_285_47# hold63/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X199 hold63/a_285_47# hold63/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X200 hold63/a_285_47# hold63/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X201 net210 hold63/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X202 VPWR acc0.A\[16\] hold74/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X203 VGND hold74/a_285_47# hold74/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X204 net221 hold74/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X205 VGND acc0.A\[16\] hold74/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X206 VPWR hold74/a_285_47# hold74/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X207 hold74/a_285_47# hold74/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X208 hold74/a_285_47# hold74/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X209 net221 hold74/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X210 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X211 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X212 VPWR _0164_ hold85/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X213 VGND hold85/a_285_47# hold85/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X214 net232 hold85/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X215 VGND _0164_ hold85/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X216 VPWR hold85/a_285_47# hold85/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X217 hold85/a_285_47# hold85/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X218 hold85/a_285_47# hold85/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X219 net232 hold85/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X220 VPWR net50 hold96/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X221 VGND hold96/a_285_47# hold96/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X222 net243 hold96/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X223 VGND net50 hold96/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X224 VPWR hold96/a_285_47# hold96/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X225 hold96/a_285_47# hold96/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X226 hold96/a_285_47# hold96/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X227 net243 hold96/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X228 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X229 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X230 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X231 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X232 _0521_/a_81_21# _0192_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08937 pd=0.925 as=0.25675 ps=1.44 w=0.65 l=0.15
X233 _0521_/a_299_297# _0192_ _0521_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.26 ps=2.52 w=1 l=0.15
X234 VPWR _0521_/a_81_21# _0151_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X235 VPWR net230 _0521_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X236 VGND _0521_/a_81_21# _0151_ VGND sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.169 ps=1.82 w=0.65 l=0.15
X237 VGND _0179_ _0521_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X238 _0521_/a_299_297# _0179_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X239 _0521_/a_384_47# net230 _0521_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08937 ps=0.925 w=0.65 l=0.15
X240 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X241 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X242 net50 _1004_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X243 _1004_/a_891_413# _1004_/a_193_47# _1004_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X244 _1004_/a_561_413# _1004_/a_27_47# _1004_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X245 VPWR net90 _1004_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X246 net50 _1004_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X247 _1004_/a_381_47# _0102_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X248 VGND _1004_/a_634_159# _1004_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X249 VPWR _1004_/a_891_413# _1004_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X250 _1004_/a_466_413# _1004_/a_193_47# _1004_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X251 VPWR _1004_/a_634_159# _1004_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X252 _1004_/a_634_159# _1004_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X253 _1004_/a_634_159# _1004_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X254 _1004_/a_975_413# _1004_/a_193_47# _1004_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X255 VGND _1004_/a_1059_315# _1004_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X256 _1004_/a_193_47# _1004_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X257 _1004_/a_891_413# _1004_/a_27_47# _1004_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X258 _1004_/a_592_47# _1004_/a_193_47# _1004_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X259 VPWR _1004_/a_1059_315# _1004_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X260 _1004_/a_1017_47# _1004_/a_27_47# _1004_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X261 _1004_/a_193_47# _1004_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X262 _1004_/a_466_413# _1004_/a_27_47# _1004_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X263 VGND _1004_/a_891_413# _1004_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X264 _1004_/a_381_47# _0102_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X265 VGND net90 _1004_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X266 VPWR _0719_/a_27_47# _0350_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X267 _0350_ _0719_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X268 VPWR control0.add _0719_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X269 _0350_ _0719_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X270 VGND _0719_/a_27_47# _0350_ VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X271 VGND control0.add _0719_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X272 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X273 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X274 VPWR output53/a_27_47# pp[25] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X275 pp[25] output53/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X276 VPWR net53 output53/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X277 pp[25] output53/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X278 VGND output53/a_27_47# pp[25] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X279 VGND net53 output53/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X280 VPWR output42/a_27_47# pp[15] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X281 pp[15] output42/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X282 VPWR net42 output42/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X283 pp[15] output42/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X284 VGND output42/a_27_47# pp[15] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X285 VGND net42 output42/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X286 VPWR net64 output64/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X287 VGND output64/a_27_47# pp[6] VGND sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X288 VGND output64/a_27_47# pp[6] VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X289 pp[6] output64/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X290 pp[6] output64/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X291 VGND net64 output64/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X292 VPWR output64/a_27_47# pp[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X293 pp[6] output64/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X294 pp[6] output64/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X295 VPWR output64/a_27_47# pp[6] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X296 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X297 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X298 VPWR _0182_ _0504_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X299 VGND _0504_/a_27_47# _0183_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X300 VGND _0504_/a_27_47# _0183_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X301 _0183_ _0504_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X302 _0183_ _0504_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X303 VGND _0182_ _0504_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X304 VPWR _0504_/a_27_47# _0183_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X305 _0183_ _0504_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X306 _0183_ _0504_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X307 VPWR _0504_/a_27_47# _0183_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X308 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X309 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X310 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X311 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X312 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X313 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X314 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X315 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X316 net58 _0984_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X317 _0984_/a_891_413# _0984_/a_193_47# _0984_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X318 _0984_/a_561_413# _0984_/a_27_47# _0984_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X319 VPWR net70 _0984_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X320 net58 _0984_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X321 _0984_/a_381_47# _0082_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X322 VGND _0984_/a_634_159# _0984_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X323 VPWR _0984_/a_891_413# _0984_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X324 _0984_/a_466_413# _0984_/a_193_47# _0984_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X325 VPWR _0984_/a_634_159# _0984_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X326 _0984_/a_634_159# _0984_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X327 _0984_/a_634_159# _0984_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X328 _0984_/a_975_413# _0984_/a_193_47# _0984_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X329 VGND _0984_/a_1059_315# _0984_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X330 _0984_/a_193_47# _0984_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X331 _0984_/a_891_413# _0984_/a_27_47# _0984_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X332 _0984_/a_592_47# _0984_/a_193_47# _0984_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X333 VPWR _0984_/a_1059_315# _0984_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X334 _0984_/a_1017_47# _0984_/a_27_47# _0984_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X335 _0984_/a_193_47# _0984_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X336 _0984_/a_466_413# _0984_/a_27_47# _0984_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X337 VGND _0984_/a_891_413# _0984_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X338 _0984_/a_381_47# _0082_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X339 VGND net70 _0984_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X340 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X341 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X342 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=2.89
X343 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=2.89
X344 _0485_ _0967_/a_215_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X345 VGND _0967_/a_215_297# _0485_ VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X346 VPWR _0967_/a_215_297# _0485_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X347 _0967_/a_109_93# control0.state\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X348 _0967_/a_215_297# _0967_/a_109_93# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.16535 ps=1.82 w=0.65 l=0.15
X349 VGND _0476_ _0967_/a_215_297# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X350 VGND control0.state\[0\] _0967_/a_215_297# VGND sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X351 _0485_ _0967_/a_215_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X352 _0967_/a_215_297# control0.state\[2\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X353 _0967_/a_109_93# control0.state\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X354 VPWR control0.state\[0\] _0967_/a_487_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X355 VGND _0967_/a_215_297# _0485_ VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X356 _0967_/a_487_297# control0.state\[2\] _0967_/a_403_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X357 _0967_/a_403_297# _0476_ _0967_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X358 VPWR _0967_/a_215_297# _0485_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X359 _0485_ _0967_/a_215_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X360 _0485_ _0967_/a_215_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X361 _0967_/a_297_297# _0967_/a_109_93# _0967_/a_215_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
X362 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X363 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X364 net139 clknet_1_0__leaf__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X365 VGND clknet_1_0__leaf__0465_ net139 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X366 net139 clknet_1_0__leaf__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X367 VPWR clknet_1_0__leaf__0465_ net139 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X368 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X369 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X370 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X371 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X372 _0752_/a_300_297# _0752_/a_27_413# _0376_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X373 VGND _0375_ _0752_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.091 ps=0.93 w=0.65 l=0.15
X374 VPWR _0234_ _0752_/a_27_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X375 _0376_ _0752_/a_27_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.10187 ps=0.99 w=0.65 l=0.15
X376 VPWR _0222_ _0752_/a_300_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X377 _0752_/a_384_47# _0222_ _0376_ VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.143 ps=1.09 w=0.65 l=0.15
X378 VGND _0234_ _0752_/a_27_413# VGND sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.1113 ps=1.37 w=0.42 l=0.15
X379 _0752_/a_300_297# _0375_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X380 VPWR _0251_ _0429_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X381 _0429_ _0251_ _0821_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X382 _0821_/a_113_47# _0252_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X383 _0429_ _0252_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X384 VPWR _0313_ _0315_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X385 _0315_ _0313_ _0683_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X386 _0683_/a_113_47# _0314_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X387 _0315_ _0314_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X388 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X389 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X390 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X391 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X392 net120 clknet_1_1__leaf__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X393 VGND clknet_1_1__leaf__0463_ net120 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X394 net120 clknet_1_1__leaf__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X395 VPWR clknet_1_1__leaf__0463_ net120 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X396 acc0.A\[20\] _1020_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X397 _1020_/a_891_413# _1020_/a_193_47# _1020_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X398 _1020_/a_561_413# _1020_/a_27_47# _1020_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X399 VPWR net106 _1020_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X400 acc0.A\[20\] _1020_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X401 _1020_/a_381_47# _0118_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X402 VGND _1020_/a_634_159# _1020_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X403 VPWR _1020_/a_891_413# _1020_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X404 _1020_/a_466_413# _1020_/a_193_47# _1020_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X405 VPWR _1020_/a_634_159# _1020_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X406 _1020_/a_634_159# _1020_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X407 _1020_/a_634_159# _1020_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X408 _1020_/a_975_413# _1020_/a_193_47# _1020_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X409 VGND _1020_/a_1059_315# _1020_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X410 _1020_/a_193_47# _1020_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X411 _1020_/a_891_413# _1020_/a_27_47# _1020_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X412 _1020_/a_592_47# _1020_/a_193_47# _1020_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X413 VPWR _1020_/a_1059_315# _1020_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X414 _1020_/a_1017_47# _1020_/a_27_47# _1020_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X415 _1020_/a_193_47# _1020_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X416 _1020_/a_466_413# _1020_/a_27_47# _1020_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X417 VGND _1020_/a_891_413# _1020_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X418 _1020_/a_381_47# _0118_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X419 VGND net106 _1020_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X420 net134 clknet_1_0__leaf__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X421 VGND clknet_1_0__leaf__0464_ net134 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X422 net134 clknet_1_0__leaf__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X423 VPWR clknet_1_0__leaf__0464_ net134 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X424 VPWR clknet_0__0458_ clkbuf_1_0__f__0458_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X425 VPWR clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X426 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X427 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X428 VPWR clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X429 VPWR clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X430 clkbuf_1_0__f__0458_/a_110_47# clknet_0__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X431 clkbuf_1_0__f__0458_/a_110_47# clknet_0__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X432 VGND clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X433 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X434 VGND clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X435 clkbuf_1_0__f__0458_/a_110_47# clknet_0__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X436 VGND clknet_0__0458_ clkbuf_1_0__f__0458_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X437 VGND clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X438 VPWR clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X439 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X440 VGND clknet_0__0458_ clkbuf_1_0__f__0458_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X441 VGND clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X442 VPWR clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X443 VGND clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X444 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X445 clkbuf_1_0__f__0458_/a_110_47# clknet_0__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X446 VPWR clknet_0__0458_ clkbuf_1_0__f__0458_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X447 VPWR clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X448 VPWR clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X449 VGND clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X450 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X451 VGND clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X452 VGND clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X453 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X454 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X455 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X456 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X457 VPWR clkbuf_1_0__f__0458_/a_110_47# clknet_1_0__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X458 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X459 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X460 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X461 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X462 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X463 clknet_1_0__leaf__0458_ clkbuf_1_0__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X464 VPWR _0350_ _0735_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X465 VGND _0350_ _0363_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X466 _0735_/a_109_297# net224 _0363_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X467 _0363_ net224 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X468 VGND _0347_ _0804_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10563 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X469 _0804_/a_510_47# _0416_ _0804_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.143 ps=1.09 w=0.65 l=0.15
X470 _0804_/a_79_21# _0399_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.175 ps=1.35 w=1 l=0.15
X471 VPWR _0416_ _0804_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.175 pd=1.35 as=0.22 ps=1.44 w=1 l=0.15
X472 _0804_/a_79_21# _0415_ _0804_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.1625 ps=1.325 w=1 l=0.15
X473 _0804_/a_297_297# _0347_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X474 _0804_/a_79_21# _0399_ _0804_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.11375 ps=1 w=0.65 l=0.15
X475 VPWR _0804_/a_79_21# _0092_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X476 VGND _0804_/a_79_21# _0092_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X477 _0804_/a_215_47# _0415_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.10563 ps=0.975 w=0.65 l=0.15
X478 VPWR acc0.A\[12\] _0298_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X479 _0298_ acc0.A\[12\] _0666_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X480 _0666_/a_113_47# net39 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X481 _0298_ net39 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X482 _0229_ _0228_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X483 VGND _0228_ _0229_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X484 _0229_ _0228_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X485 VPWR _0228_ _0229_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X486 VPWR control0.count\[3\] hold20/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X487 VGND hold20/a_285_47# hold20/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X488 net167 hold20/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X489 VGND control0.count\[3\] hold20/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X490 VPWR hold20/a_285_47# hold20/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X491 hold20/a_285_47# hold20/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X492 hold20/a_285_47# hold20/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X493 net167 hold20/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X494 VPWR acc0.A\[8\] hold31/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X495 VGND hold31/a_285_47# hold31/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X496 net178 hold31/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X497 VGND acc0.A\[8\] hold31/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X498 VPWR hold31/a_285_47# hold31/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X499 hold31/a_285_47# hold31/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X500 hold31/a_285_47# hold31/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X501 net178 hold31/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X502 VPWR _0155_ hold42/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X503 VGND hold42/a_285_47# hold42/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X504 net189 hold42/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X505 VGND _0155_ hold42/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X506 VPWR hold42/a_285_47# hold42/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X507 hold42/a_285_47# hold42/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X508 hold42/a_285_47# hold42/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X509 net189 hold42/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X510 VPWR _0123_ hold53/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X511 VGND hold53/a_285_47# hold53/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X512 net200 hold53/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X513 VGND _0123_ hold53/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X514 VPWR hold53/a_285_47# hold53/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X515 hold53/a_285_47# hold53/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X516 hold53/a_285_47# hold53/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X517 net200 hold53/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X518 VPWR acc0.A\[19\] hold64/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X519 VGND hold64/a_285_47# hold64/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X520 net211 hold64/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X521 VGND acc0.A\[19\] hold64/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X522 VPWR hold64/a_285_47# hold64/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X523 hold64/a_285_47# hold64/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X524 hold64/a_285_47# hold64/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X525 net211 hold64/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X526 VPWR net58 hold75/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X527 VGND hold75/a_285_47# hold75/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X528 net222 hold75/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X529 VGND net58 hold75/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X530 VPWR hold75/a_285_47# hold75/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X531 hold75/a_285_47# hold75/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X532 hold75/a_285_47# hold75/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X533 net222 hold75/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X534 VPWR net61 hold86/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X535 VGND hold86/a_285_47# hold86/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X536 net233 hold86/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X537 VGND net61 hold86/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X538 VPWR hold86/a_285_47# hold86/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X539 hold86/a_285_47# hold86/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X540 hold86/a_285_47# hold86/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X541 net233 hold86/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X542 VPWR net54 hold97/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X543 VGND hold97/a_285_47# hold97/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X544 net244 hold97/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X545 VGND net54 hold97/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X546 VPWR hold97/a_285_47# hold97/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X547 hold97/a_285_47# hold97/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X548 hold97/a_285_47# hold97/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X549 net244 hold97/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X550 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X551 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X552 VPWR net14 _0520_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.16 ps=1.32 w=1 l=0.15
X553 _0520_/a_27_297# _0186_ _0520_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X554 VGND net14 _0520_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.11375 ps=1 w=0.65 l=0.15
X555 _0192_ _0520_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.155 ps=1.31 w=1 l=0.15
X556 _0520_/a_27_297# _0186_ _0520_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.25285 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X557 _0520_/a_109_297# _0180_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.2529 ps=2.52 w=1 l=0.15
X558 _0520_/a_373_47# _0180_ _0520_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.169 ps=1.82 w=0.65 l=0.15
X559 _0192_ _0520_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10075 ps=0.96 w=0.65 l=0.15
X560 _0520_/a_109_297# net168 _0520_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X561 _0520_/a_109_47# net168 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X562 net49 _1003_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X563 _1003_/a_891_413# _1003_/a_193_47# _1003_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X564 _1003_/a_561_413# _1003_/a_27_47# _1003_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X565 VPWR net89 _1003_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X566 net49 _1003_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X567 _1003_/a_381_47# _0101_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X568 VGND _1003_/a_634_159# _1003_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X569 VPWR _1003_/a_891_413# _1003_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X570 _1003_/a_466_413# _1003_/a_193_47# _1003_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X571 VPWR _1003_/a_634_159# _1003_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X572 _1003_/a_634_159# _1003_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X573 _1003_/a_634_159# _1003_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X574 _1003_/a_975_413# _1003_/a_193_47# _1003_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X575 VGND _1003_/a_1059_315# _1003_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X576 _1003_/a_193_47# _1003_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X577 _1003_/a_891_413# _1003_/a_27_47# _1003_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X578 _1003_/a_592_47# _1003_/a_193_47# _1003_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X579 VPWR _1003_/a_1059_315# _1003_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X580 _1003_/a_1017_47# _1003_/a_27_47# _1003_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X581 _1003_/a_193_47# _1003_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X582 _1003_/a_466_413# _1003_/a_27_47# _1003_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X583 VGND _1003_/a_891_413# _1003_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X584 _1003_/a_381_47# _0101_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X585 VGND net89 _1003_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X586 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X587 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X588 _0718_/a_377_297# _0337_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.365 ps=1.73 w=1 l=0.15
X589 _0718_/a_47_47# _0348_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X590 _0718_/a_129_47# _0348_ _0718_/a_47_47# VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X591 _0718_/a_285_47# _0348_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X592 _0349_ _0718_/a_47_47# _0718_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.08775 ps=0.92 w=0.65 l=0.15
X593 VGND _0337_ _0718_/a_129_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.06825 ps=0.86 w=0.65 l=0.15
X594 VPWR _0337_ _0718_/a_47_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.365 pd=1.73 as=0.135 ps=1.27 w=1 l=0.15
X595 VPWR _0718_/a_47_47# _0349_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.165 ps=1.33 w=1 l=0.15
X596 _0349_ _0348_ _0718_/a_377_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X597 _0718_/a_285_47# _0337_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X598 VPWR acc0.A\[10\] _0281_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X599 _0281_ acc0.A\[10\] _0649_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X600 _0649_/a_113_47# net37 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X601 _0281_ net37 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X602 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X603 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X604 net115 clknet_1_1__leaf__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X605 VGND clknet_1_1__leaf__0462_ net115 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X606 net115 clknet_1_1__leaf__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X607 VPWR clknet_1_1__leaf__0462_ net115 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X608 VPWR output54/a_27_47# pp[26] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X609 pp[26] output54/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X610 VPWR net54 output54/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X611 pp[26] output54/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X612 VGND output54/a_27_47# pp[26] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X613 VGND net54 output54/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X614 VPWR output43/a_27_47# pp[16] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X615 pp[16] output43/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X616 VPWR net43 output43/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X617 pp[16] output43/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X618 VGND output43/a_27_47# pp[16] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X619 VGND net43 output43/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X620 VPWR net65 output65/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X621 VGND output65/a_27_47# pp[7] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X622 VGND output65/a_27_47# pp[7] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X623 pp[7] output65/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X624 pp[7] output65/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X625 VGND net65 output65/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X626 VPWR output65/a_27_47# pp[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X627 pp[7] output65/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X628 pp[7] output65/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X629 VPWR output65/a_27_47# pp[7] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X630 VPWR _0180_ _0503_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X631 VGND _0180_ _0182_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X632 _0503_/a_109_297# control0.sh _0182_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X633 _0182_ control0.sh VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X634 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X635 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X636 net47 _0983_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X637 _0983_/a_891_413# _0983_/a_193_47# _0983_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X638 _0983_/a_561_413# _0983_/a_27_47# _0983_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X639 VPWR net69 _0983_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X640 net47 _0983_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X641 _0983_/a_381_47# _0081_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X642 VGND _0983_/a_634_159# _0983_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X643 VPWR _0983_/a_891_413# _0983_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X644 _0983_/a_466_413# _0983_/a_193_47# _0983_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X645 VPWR _0983_/a_634_159# _0983_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X646 _0983_/a_634_159# _0983_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X647 _0983_/a_634_159# _0983_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X648 _0983_/a_975_413# _0983_/a_193_47# _0983_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X649 VGND _0983_/a_1059_315# _0983_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X650 _0983_/a_193_47# _0983_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X651 _0983_/a_891_413# _0983_/a_27_47# _0983_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X652 _0983_/a_592_47# _0983_/a_193_47# _0983_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X653 VPWR _0983_/a_1059_315# _0983_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X654 _0983_/a_1017_47# _0983_/a_27_47# _0983_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X655 _0983_/a_193_47# _0983_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X656 _0983_/a_466_413# _0983_/a_27_47# _0983_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X657 VGND _0983_/a_891_413# _0983_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X658 _0983_/a_381_47# _0081_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X659 VGND net69 _0983_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X660 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X661 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X662 _0484_ _0483_ _0966_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X663 VPWR net236 _0484_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.182 pd=1.92 as=0.174 ps=1.39 w=0.7 l=0.15
X664 _0966_/a_27_47# _0483_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X665 _0484_ net236 _0966_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X666 _0966_/a_109_297# _0482_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X667 VGND _0482_ _0966_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X668 _0375_ _0751_/a_29_53# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X669 _0751_/a_111_297# _0374_ _0751_/a_29_53# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X670 _0375_ _0751_/a_29_53# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.10187 ps=0.99 w=0.65 l=0.15
X671 _0751_/a_183_297# _0227_ _0751_/a_111_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X672 VPWR _0225_ _0751_/a_183_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X673 _0751_/a_29_53# _0227_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X674 VGND _0374_ _0751_/a_29_53# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X675 VGND _0225_ _0751_/a_29_53# VGND sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X676 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X677 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X678 VGND _0369_ _0820_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X679 _0820_/a_510_47# _0428_ _0820_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X680 _0820_/a_79_21# _0399_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X681 VPWR _0428_ _0820_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X682 _0820_/a_79_21# net214 _0820_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X683 _0820_/a_297_297# _0369_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X684 _0820_/a_79_21# _0399_ _0820_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X685 VPWR _0820_/a_79_21# _0088_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X686 VGND _0820_/a_79_21# _0088_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X687 _0820_/a_215_47# net214 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X688 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X689 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X690 VGND acc0.A\[25\] _0682_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X691 _0682_/a_68_297# net53 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X692 _0314_ _0682_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X693 VPWR acc0.A\[25\] _0682_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X694 _0314_ _0682_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X695 _0682_/a_150_297# net53 _0682_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X696 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X697 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X698 VPWR _0468_ _0949_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X699 _0469_ _0949_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X700 VGND _0468_ _0949_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X701 _0949_/a_59_75# control0.state\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X702 _0469_ _0949_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X703 _0949_/a_145_75# control0.state\[0\] _0949_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X704 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X705 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X706 VGND _0218_ _0803_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X707 _0803_/a_68_297# net39 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X708 _0416_ _0803_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X709 VPWR _0218_ _0803_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X710 _0416_ _0803_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X711 _0803_/a_150_297# net39 _0803_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X712 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X713 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X714 VPWR clknet_0__0457_ clkbuf_1_0__f__0457_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X715 VPWR clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X716 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X717 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X718 VPWR clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X719 VPWR clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X720 clkbuf_1_0__f__0457_/a_110_47# clknet_0__0457_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X721 clkbuf_1_0__f__0457_/a_110_47# clknet_0__0457_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X722 VGND clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X723 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X724 VGND clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X725 clkbuf_1_0__f__0457_/a_110_47# clknet_0__0457_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X726 VGND clknet_0__0457_ clkbuf_1_0__f__0457_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X727 VGND clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X728 VPWR clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X729 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X730 VGND clknet_0__0457_ clkbuf_1_0__f__0457_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X731 VGND clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X732 VPWR clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X733 VGND clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X734 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X735 clkbuf_1_0__f__0457_/a_110_47# clknet_0__0457_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X736 VPWR clknet_0__0457_ clkbuf_1_0__f__0457_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X737 VPWR clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X738 VPWR clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X739 VGND clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X740 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X741 VGND clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X742 VGND clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X743 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X744 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X745 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X746 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X747 VPWR clkbuf_1_0__f__0457_/a_110_47# clknet_1_0__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X748 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X749 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X750 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X751 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X752 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X753 clknet_1_0__leaf__0457_ clkbuf_1_0__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X754 VPWR acc0.A\[13\] _0665_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X755 VGND acc0.A\[13\] _0297_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X756 _0665_/a_109_297# net40 _0297_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X757 _0297_ net40 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X758 _0734_/a_377_297# _0318_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=2.42 as=0 ps=0 w=1 l=0.15
X759 _0734_/a_47_47# _0361_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X760 _0734_/a_129_47# _0361_ _0734_/a_47_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.72 as=0.169 ps=1.82 w=0.65 l=0.15
X761 _0734_/a_285_47# _0361_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X762 _0362_ _0734_/a_47_47# _0734_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X763 VGND _0318_ _0734_/a_129_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X764 VPWR _0318_ _0734_/a_47_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X765 VPWR _0734_/a_47_47# _0362_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.33 ps=2.66 w=1 l=0.15
X766 _0362_ _0361_ _0734_/a_377_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X767 _0734_/a_285_47# _0318_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X768 VPWR net49 _0596_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X769 _0228_ _0596_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X770 VGND net49 _0596_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X771 _0596_/a_59_75# acc0.A\[21\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X772 _0228_ _0596_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X773 _0596_/a_145_75# acc0.A\[21\] _0596_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X774 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X775 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X776 VPWR comp0.B\[15\] hold10/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X777 VGND hold10/a_285_47# hold10/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X778 net157 hold10/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X779 VGND comp0.B\[15\] hold10/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X780 VPWR hold10/a_285_47# hold10/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X781 hold10/a_285_47# hold10/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X782 hold10/a_285_47# hold10/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X783 net157 hold10/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X784 VPWR acc0.A\[7\] hold21/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X785 VGND hold21/a_285_47# hold21/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X786 net168 hold21/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X787 VGND acc0.A\[7\] hold21/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X788 VPWR hold21/a_285_47# hold21/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X789 hold21/a_285_47# hold21/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X790 hold21/a_285_47# hold21/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X791 net168 hold21/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X792 VPWR _0153_ hold32/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X793 VGND hold32/a_285_47# hold32/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X794 net179 hold32/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X795 VGND _0153_ hold32/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X796 VPWR hold32/a_285_47# hold32/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X797 hold32/a_285_47# hold32/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X798 hold32/a_285_47# hold32/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X799 net179 hold32/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X800 VPWR acc0.A\[28\] hold43/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X801 VGND hold43/a_285_47# hold43/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X802 net190 hold43/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X803 VGND acc0.A\[28\] hold43/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X804 VPWR hold43/a_285_47# hold43/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X805 hold43/a_285_47# hold43/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X806 hold43/a_285_47# hold43/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X807 net190 hold43/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X808 VPWR comp0.B\[1\] hold54/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X809 VGND hold54/a_285_47# hold54/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X810 net201 hold54/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X811 VGND comp0.B\[1\] hold54/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X812 VPWR hold54/a_285_47# hold54/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X813 hold54/a_285_47# hold54/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X814 hold54/a_285_47# hold54/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X815 net201 hold54/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X816 VPWR net65 hold65/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X817 VGND hold65/a_285_47# hold65/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X818 net212 hold65/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X819 VGND net65 hold65/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X820 VPWR hold65/a_285_47# hold65/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X821 hold65/a_285_47# hold65/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X822 hold65/a_285_47# hold65/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X823 net212 hold65/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X824 VPWR net46 hold76/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X825 VGND hold76/a_285_47# hold76/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X826 net223 hold76/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X827 VGND net46 hold76/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X828 VPWR hold76/a_285_47# hold76/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X829 hold76/a_285_47# hold76/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X830 hold76/a_285_47# hold76/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X831 net223 hold76/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X832 VPWR net36 hold87/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X833 VGND hold87/a_285_47# hold87/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X834 net234 hold87/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X835 VGND net36 hold87/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X836 VPWR hold87/a_285_47# hold87/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X837 hold87/a_285_47# hold87/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X838 hold87/a_285_47# hold87/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X839 net234 hold87/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X840 VPWR net40 hold98/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X841 VGND hold98/a_285_47# hold98/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X842 net245 hold98/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X843 VGND net40 hold98/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X844 VPWR hold98/a_285_47# hold98/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X845 hold98/a_285_47# hold98/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X846 hold98/a_285_47# hold98/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X847 net245 hold98/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X848 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X849 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X850 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X851 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X852 net48 _1002_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X853 _1002_/a_891_413# _1002_/a_193_47# _1002_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X854 _1002_/a_561_413# _1002_/a_27_47# _1002_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X855 VPWR net88 _1002_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X856 net48 _1002_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X857 _1002_/a_381_47# _0100_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X858 VGND _1002_/a_634_159# _1002_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X859 VPWR _1002_/a_891_413# _1002_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X860 _1002_/a_466_413# _1002_/a_193_47# _1002_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X861 VPWR _1002_/a_634_159# _1002_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X862 _1002_/a_634_159# _1002_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X863 _1002_/a_634_159# _1002_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X864 _1002_/a_975_413# _1002_/a_193_47# _1002_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X865 VGND _1002_/a_1059_315# _1002_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X866 _1002_/a_193_47# _1002_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X867 _1002_/a_891_413# _1002_/a_27_47# _1002_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X868 _1002_/a_592_47# _1002_/a_193_47# _1002_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X869 VPWR _1002_/a_1059_315# _1002_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X870 _1002_/a_1017_47# _1002_/a_27_47# _1002_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X871 _1002_/a_193_47# _1002_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X872 _1002_/a_466_413# _1002_/a_27_47# _1002_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X873 VGND _1002_/a_891_413# _1002_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X874 _1002_/a_381_47# _0100_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X875 VGND net88 _1002_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X876 _0648_/a_27_297# _0277_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X877 _0648_/a_27_297# _0279_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X878 _0648_/a_277_297# _0277_ _0648_/a_205_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X879 VPWR _0276_ _0648_/a_277_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X880 _0280_ _0648_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.10187 ps=0.99 w=0.65 l=0.15
X881 _0648_/a_205_297# _0278_ _0648_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X882 _0280_ _0648_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X883 VGND _0278_ _0648_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X884 _0648_/a_109_297# _0279_ _0648_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X885 VGND _0276_ _0648_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X886 VPWR _0717_/a_80_21# _0348_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X887 _0717_/a_209_297# _0334_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X888 _0717_/a_303_47# _0333_ _0717_/a_209_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X889 _0717_/a_209_47# _0334_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.11213 ps=0.995 w=0.65 l=0.15
X890 VGND _0717_/a_80_21# _0348_ VGND sky130_fd_pr__nfet_01v8 ad=0.11213 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X891 VGND _0335_ _0717_/a_80_21# VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X892 _0717_/a_80_21# _0221_ _0717_/a_303_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X893 VPWR _0333_ _0717_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X894 _0717_/a_80_21# _0335_ _0717_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X895 _0717_/a_209_297# _0221_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
X896 VPWR _0183_ _0579_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X897 _0579_/a_27_297# _0217_ _0579_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X898 VGND _0183_ _0579_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X899 _0118_ _0579_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X900 _0579_/a_27_297# _0217_ _0579_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X901 _0579_/a_109_297# net187 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X902 _0579_/a_373_47# net187 _0579_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X903 _0118_ _0579_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X904 _0579_/a_109_297# net211 _0579_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X905 _0579_/a_109_47# net211 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X906 VPWR output55/a_27_47# pp[27] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X907 pp[27] output55/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X908 VPWR net55 output55/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X909 pp[27] output55/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X910 VGND output55/a_27_47# pp[27] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X911 VGND net55 output55/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X912 VPWR output44/a_27_47# pp[17] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X913 pp[17] output44/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X914 VPWR net44 output44/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X915 pp[17] output44/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X916 VGND output44/a_27_47# pp[17] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X917 VGND net44 output44/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X918 VPWR net66 output66/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X919 VGND output66/a_27_47# pp[8] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X920 VGND output66/a_27_47# pp[8] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X921 pp[8] output66/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X922 pp[8] output66/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X923 VGND net66 output66/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X924 VPWR output66/a_27_47# pp[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X925 pp[8] output66/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X926 pp[8] output66/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X927 VPWR output66/a_27_47# pp[8] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X928 net68 clknet_1_0__leaf__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X929 VGND clknet_1_0__leaf__0458_ net68 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X930 net68 clknet_1_0__leaf__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X931 VPWR clknet_1_0__leaf__0458_ net68 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X932 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X933 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X934 VPWR _0180_ _0502_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X935 VGND _0502_/a_27_47# _0181_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X936 VGND _0502_/a_27_47# _0181_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X937 _0181_ _0502_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X938 _0181_ _0502_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X939 VGND _0180_ _0502_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X940 VPWR _0502_/a_27_47# _0181_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X941 _0181_ _0502_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X942 _0181_ _0502_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X943 VPWR _0502_/a_27_47# _0181_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X944 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X945 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X946 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X947 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X948 net93 clknet_1_1__leaf__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X949 VGND clknet_1_1__leaf__0460_ net93 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X950 net93 clknet_1_1__leaf__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X951 VPWR clknet_1_1__leaf__0460_ net93 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X952 net36 _0982_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X953 _0982_/a_891_413# _0982_/a_193_47# _0982_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X954 _0982_/a_561_413# _0982_/a_27_47# _0982_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X955 VPWR net68 _0982_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X956 net36 _0982_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X957 _0982_/a_381_47# _0080_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X958 VGND _0982_/a_634_159# _0982_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X959 VPWR _0982_/a_891_413# _0982_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X960 _0982_/a_466_413# _0982_/a_193_47# _0982_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X961 VPWR _0982_/a_634_159# _0982_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X962 _0982_/a_634_159# _0982_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X963 _0982_/a_634_159# _0982_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X964 _0982_/a_975_413# _0982_/a_193_47# _0982_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X965 VGND _0982_/a_1059_315# _0982_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X966 _0982_/a_193_47# _0982_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X967 _0982_/a_891_413# _0982_/a_27_47# _0982_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X968 _0982_/a_592_47# _0982_/a_193_47# _0982_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X969 VPWR _0982_/a_1059_315# _0982_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X970 _0982_/a_1017_47# _0982_/a_27_47# _0982_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X971 _0982_/a_193_47# _0982_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X972 _0982_/a_466_413# _0982_/a_27_47# _0982_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X973 VGND _0982_/a_891_413# _0982_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X974 _0982_/a_381_47# _0080_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X975 VGND net68 _0982_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X976 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X977 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X978 _0965_/a_377_297# control0.count\[3\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=2.42 as=0 ps=0 w=1 l=0.15
X979 _0965_/a_47_47# _0478_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X980 _0965_/a_129_47# _0478_ _0965_/a_47_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.72 as=0.169 ps=1.82 w=0.65 l=0.15
X981 _0965_/a_285_47# _0478_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X982 _0483_ _0965_/a_47_47# _0965_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X983 VGND control0.count\[3\] _0965_/a_129_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X984 VPWR control0.count\[3\] _0965_/a_47_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X985 VPWR _0965_/a_47_47# _0483_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.33 ps=2.66 w=1 l=0.15
X986 _0483_ _0478_ _0965_/a_377_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X987 _0965_/a_285_47# control0.count\[3\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X988 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X989 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X990 VPWR acc0.A\[25\] _0313_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X991 _0313_ acc0.A\[25\] _0681_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X992 _0681_/a_113_47# net53 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X993 _0313_ net53 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X994 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X995 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X996 VPWR _0226_ _0750_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2415 ps=2.83 w=0.42 l=0.15
X997 VPWR _0373_ _0750_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X998 _0750_/a_181_47# _0229_ _0750_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0882 pd=1.26 as=0.0882 ps=1.26 w=0.42 l=0.15
X999 VGND _0373_ _0750_/a_181_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1000 _0750_/a_27_47# _0229_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1001 _0374_ _0750_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1002 _0374_ _0750_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1003 _0750_/a_109_47# _0226_ _0750_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1004 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1005 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1006 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X1007 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X1008 VPWR net34 _0948_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X1009 VGND net34 _0468_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1010 _0948_/a_109_297# control0.state\[2\] _0468_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1011 _0468_ control0.state\[2\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1012 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1013 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1014 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1015 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1016 VPWR _0414_ _0802_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X1017 _0415_ _0802_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X1018 VGND _0414_ _0802_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X1019 _0802_/a_59_75# _0404_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1020 _0415_ _0802_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X1021 _0802_/a_145_75# _0404_ _0802_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X1022 VPWR _0281_ _0664_/a_382_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.305 ps=2.61 w=1 l=0.15
X1023 _0664_/a_297_47# _0285_ _0664_/a_79_21# VGND sky130_fd_pr__nfet_01v8 ad=0.3705 pd=3.74 as=0.169 ps=1.82 w=0.65 l=0.15
X1024 _0664_/a_297_47# _0281_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1025 VGND _0284_ _0664_/a_297_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1026 VPWR _0664_/a_79_21# _0296_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.28 ps=2.56 w=1 l=0.15
X1027 _0664_/a_79_21# _0285_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.15
X1028 _0664_/a_382_297# _0284_ _0664_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1029 VGND _0664_/a_79_21# _0296_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1030 _0733_/a_222_93# _0319_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X1031 VPWR _0321_ _0733_/a_544_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X1032 VGND _0733_/a_79_199# _0361_ VGND sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X1033 _0733_/a_222_93# _0319_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.18575 ps=1.415 w=0.42 l=0.15
X1034 VGND _0360_ _0733_/a_448_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1035 _0733_/a_448_47# _0733_/a_222_93# _0733_/a_79_199# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X1036 _0733_/a_79_199# _0733_/a_222_93# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X1037 _0733_/a_544_297# _0360_ _0733_/a_79_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X1038 _0733_/a_448_47# _0321_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X1039 VPWR _0733_/a_79_199# _0361_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18575 pd=1.415 as=0.26 ps=2.52 w=1 l=0.15
X1040 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1041 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1042 VPWR acc0.A\[21\] _0595_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X1043 VGND acc0.A\[21\] _0227_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1044 _0595_/a_109_297# net49 _0227_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1045 _0227_ net49 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1046 VPWR _0144_ hold11/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1047 VGND hold11/a_285_47# hold11/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1048 net158 hold11/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1049 VGND _0144_ hold11/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1050 VPWR hold11/a_285_47# hold11/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1051 hold11/a_285_47# hold11/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1052 hold11/a_285_47# hold11/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1053 net158 hold11/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1054 VPWR _0152_ hold22/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1055 VGND hold22/a_285_47# hold22/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1056 net169 hold22/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1057 VGND _0152_ hold22/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1058 VPWR hold22/a_285_47# hold22/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1059 hold22/a_285_47# hold22/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1060 hold22/a_285_47# hold22/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1061 net169 hold22/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1062 VPWR comp0.B\[8\] hold33/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1063 VGND hold33/a_285_47# hold33/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1064 net180 hold33/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1065 VGND comp0.B\[8\] hold33/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1066 VPWR hold33/a_285_47# hold33/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1067 hold33/a_285_47# hold33/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1068 hold33/a_285_47# hold33/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1069 net180 hold33/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1070 VPWR _0127_ hold44/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1071 VGND hold44/a_285_47# hold44/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1072 net191 hold44/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1073 VGND _0127_ hold44/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1074 VPWR hold44/a_285_47# hold44/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1075 hold44/a_285_47# hold44/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1076 hold44/a_285_47# hold44/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1077 net191 hold44/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1078 VPWR _0130_ hold55/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1079 VGND hold55/a_285_47# hold55/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1080 net202 hold55/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1081 VGND _0130_ hold55/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1082 VPWR hold55/a_285_47# hold55/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1083 hold55/a_285_47# hold55/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1084 hold55/a_285_47# hold55/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1085 net202 hold55/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1086 VPWR net49 hold66/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1087 VGND hold66/a_285_47# hold66/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1088 net213 hold66/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1089 VGND net49 hold66/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1090 VPWR hold66/a_285_47# hold66/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1091 hold66/a_285_47# hold66/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1092 hold66/a_285_47# hold66/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1093 net213 hold66/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1094 VPWR net55 hold77/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1095 VGND hold77/a_285_47# hold77/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1096 net224 hold77/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1097 VGND net55 hold77/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1098 VPWR hold77/a_285_47# hold77/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1099 hold77/a_285_47# hold77/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1100 hold77/a_285_47# hold77/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1101 net224 hold77/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1102 VPWR net64 hold88/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1103 VGND hold88/a_285_47# hold88/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1104 net235 hold88/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1105 VGND net64 hold88/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1106 VPWR hold88/a_285_47# hold88/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1107 hold88/a_285_47# hold88/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1108 hold88/a_285_47# hold88/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1109 net235 hold88/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1110 VPWR net38 hold99/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1111 VGND hold99/a_285_47# hold99/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1112 net246 hold99/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1113 VGND net38 hold99/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1114 VPWR hold99/a_285_47# hold99/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1115 hold99/a_285_47# hold99/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1116 hold99/a_285_47# hold99/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1117 net246 hold99/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1118 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1119 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1120 net46 _1001_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1121 _1001_/a_891_413# _1001_/a_193_47# _1001_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X1122 _1001_/a_561_413# _1001_/a_27_47# _1001_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X1123 VPWR net87 _1001_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1124 net46 _1001_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1125 _1001_/a_381_47# _0099_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X1126 VGND _1001_/a_634_159# _1001_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X1127 VPWR _1001_/a_891_413# _1001_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1128 _1001_/a_466_413# _1001_/a_193_47# _1001_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1129 VPWR _1001_/a_634_159# _1001_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1130 _1001_/a_634_159# _1001_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X1131 _1001_/a_634_159# _1001_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X1132 _1001_/a_975_413# _1001_/a_193_47# _1001_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X1133 VGND _1001_/a_1059_315# _1001_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X1134 _1001_/a_193_47# _1001_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X1135 _1001_/a_891_413# _1001_/a_27_47# _1001_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1136 _1001_/a_592_47# _1001_/a_193_47# _1001_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X1137 VPWR _1001_/a_1059_315# _1001_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1138 _1001_/a_1017_47# _1001_/a_27_47# _1001_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X1139 _1001_/a_193_47# _1001_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X1140 _1001_/a_466_413# _1001_/a_27_47# _1001_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X1141 VGND _1001_/a_891_413# _1001_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1142 _1001_/a_381_47# _0099_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1143 VGND net87 _1001_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1144 VPWR _0346_ _0716_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X1145 VGND _0716_/a_27_47# _0347_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X1146 VGND _0716_/a_27_47# _0347_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1147 _0347_ _0716_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X1148 _0347_ _0716_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1149 VGND _0346_ _0716_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X1150 VPWR _0716_/a_27_47# _0347_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1151 _0347_ _0716_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1152 _0347_ _0716_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1153 VPWR _0716_/a_27_47# _0347_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1154 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1155 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1156 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1157 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1158 VPWR _0183_ _0578_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X1159 _0578_/a_27_297# _0217_ _0578_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X1160 VGND _0183_ _0578_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X1161 _0119_ _0578_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1162 _0578_/a_27_297# _0217_ _0578_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X1163 _0578_/a_109_297# net150 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1164 _0578_/a_373_47# net150 _0578_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1165 _0119_ _0578_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1166 _0578_/a_109_297# net187 _0578_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1167 _0578_/a_109_47# net187 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1168 _0647_/a_377_297# acc0.A\[12\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=2.42 as=0 ps=0 w=1 l=0.15
X1169 _0647_/a_47_47# net39 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1170 _0647_/a_129_47# net39 _0647_/a_47_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.72 as=0.169 ps=1.82 w=0.65 l=0.15
X1171 _0647_/a_285_47# net39 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X1172 _0279_ _0647_/a_47_47# _0647_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X1173 VGND acc0.A\[12\] _0647_/a_129_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1174 VPWR acc0.A\[12\] _0647_/a_47_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1175 VPWR _0647_/a_47_47# _0279_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.33 ps=2.66 w=1 l=0.15
X1176 _0279_ net39 _0647_/a_377_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1177 _0647_/a_285_47# acc0.A\[12\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1178 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1179 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1180 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1181 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1182 VPWR output56/a_27_47# pp[28] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1183 pp[28] output56/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1184 VPWR net56 output56/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1185 pp[28] output56/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X1186 VGND output56/a_27_47# pp[28] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1187 VGND net56 output56/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1188 VPWR output45/a_27_47# pp[18] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1189 pp[18] output45/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1190 VPWR net45 output45/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1191 pp[18] output45/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X1192 VGND output45/a_27_47# pp[18] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1193 VGND net45 output45/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1194 VPWR net67 output67/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X1195 VGND output67/a_27_47# pp[9] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X1196 VGND output67/a_27_47# pp[9] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1197 pp[9] output67/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X1198 pp[9] output67/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1199 VGND net67 output67/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X1200 VPWR output67/a_27_47# pp[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1201 pp[9] output67/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1202 pp[9] output67/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1203 VPWR output67/a_27_47# pp[9] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1204 VPWR _0501_/a_27_47# _0180_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1205 _0180_ _0501_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1206 VPWR control0.reset _0501_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1207 _0180_ _0501_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X1208 VGND _0501_/a_27_47# _0180_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1209 VGND control0.reset _0501_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1210 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X1211 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X1212 net70 clknet_1_0__leaf__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1213 VGND clknet_1_0__leaf__0458_ net70 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1214 net70 clknet_1_0__leaf__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1215 VPWR clknet_1_0__leaf__0458_ net70 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1216 VPWR _0466_ _0981_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X1217 _0981_/a_27_297# _0490_ _0981_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X1218 VGND _0466_ _0981_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X1219 _0170_ _0981_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1220 _0981_/a_27_297# _0490_ _0981_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X1221 _0981_/a_109_297# net167 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1222 _0981_/a_373_47# net167 _0981_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1223 _0170_ _0981_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1224 _0981_/a_109_297# _0488_ _0981_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1225 _0981_/a_109_47# _0488_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1226 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X1227 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X1228 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1229 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1230 VPWR _0480_ _0964_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X1231 VGND _0480_ _0482_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1232 _0964_/a_109_297# _0481_ _0482_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1233 _0482_ _0481_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1234 net131 clknet_1_1__leaf__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1235 VGND clknet_1_1__leaf__0464_ net131 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1236 net131 clknet_1_1__leaf__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1237 VPWR clknet_1_1__leaf__0464_ net131 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1238 net145 clknet_1_1__leaf__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1239 VGND clknet_1_1__leaf__0465_ net145 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1240 net145 clknet_1_1__leaf__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1241 VPWR clknet_1_1__leaf__0465_ net145 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1242 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1243 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1244 VPWR _0680_/a_80_21# _0312_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.265 ps=2.53 w=1 l=0.15
X1245 _0680_/a_80_21# _0238_ _0680_/a_472_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.155 ps=1.31 w=1 l=0.15
X1246 VPWR _0305_ _0680_/a_217_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1247 VGND _0311_ _0680_/a_80_21# VGND sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.091 ps=0.93 w=0.65 l=0.15
X1248 VGND _0680_/a_80_21# _0312_ VGND sky130_fd_pr__nfet_01v8 ad=0.26 pd=1.45 as=0.17225 ps=1.83 w=0.65 l=0.15
X1249 _0680_/a_300_47# _0305_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.26 ps=1.45 w=0.65 l=0.15
X1250 _0680_/a_217_297# _0294_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1251 _0680_/a_80_21# _0294_ _0680_/a_300_47# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.091 ps=0.93 w=0.65 l=0.15
X1252 _0680_/a_472_297# _0311_ _0680_/a_217_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.155 pd=1.31 as=0.14 ps=1.28 w=1 l=0.15
X1253 _0680_/a_80_21# _0238_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.10075 ps=0.96 w=0.65 l=0.15
X1254 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1255 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1256 net78 clknet_1_1__leaf__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1257 VGND clknet_1_1__leaf__0459_ net78 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1258 net78 clknet_1_1__leaf__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1259 VPWR clknet_1_1__leaf__0459_ net78 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1260 VPWR control0.state\[2\] _0947_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X1261 VGND control0.state\[2\] _0467_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1262 _0947_/a_109_297# _0466_ _0467_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1263 _0467_ _0466_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1264 VPWR clknet_1_0__leaf_clk clkload0/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X1265 VGND clkload0/a_27_47# clkload0/X VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X1266 VGND clkload0/a_27_47# clkload0/X VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1267 clkload0/X clkload0/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X1268 clkload0/X clkload0/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1269 VGND clknet_1_0__leaf_clk clkload0/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X1270 VPWR clkload0/a_27_47# clkload0/X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1271 clkload0/X clkload0/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1272 clkload0/X clkload0/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1273 VPWR clkload0/a_27_47# clkload0/X VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1274 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1275 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1276 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1277 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1278 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1279 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1280 VPWR _0279_ _0414_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1281 _0414_ _0279_ _0801_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X1282 _0801_/a_113_47# _0403_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1283 _0414_ _0403_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1284 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1285 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1286 VPWR _0290_ _0663_/a_207_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1287 _0295_ _0663_/a_207_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X1288 _0663_/a_297_47# _0663_/a_27_413# _0663_/a_207_413# VGND sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X1289 _0295_ _0663_/a_207_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X1290 _0663_/a_207_413# _0663_/a_27_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X1291 VPWR _0288_ _0663_/a_27_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X1292 VGND _0290_ _0663_/a_297_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X1293 _0663_/a_27_413# _0288_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1294 VPWR _0732_/a_80_21# _0360_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X1295 _0732_/a_209_297# _0313_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.65 pd=5.3 as=0 ps=0 w=1 l=0.15
X1296 _0732_/a_303_47# _0359_ _0732_/a_209_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.208 ps=1.94 w=0.65 l=0.15
X1297 _0732_/a_209_47# _0313_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1298 VGND _0732_/a_80_21# _0360_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.17225 ps=1.83 w=0.65 l=0.15
X1299 VGND _0328_ _0732_/a_80_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2145 ps=1.96 w=0.65 l=0.15
X1300 _0732_/a_80_21# _0324_ _0732_/a_303_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1301 VPWR _0359_ _0732_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1302 _0732_/a_80_21# _0328_ _0732_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0 ps=0 w=1 l=0.15
X1303 _0732_/a_209_297# _0324_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1304 VPWR acc0.A\[20\] _0226_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1305 _0226_ acc0.A\[20\] _0594_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X1306 _0594_/a_113_47# net48 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1307 _0226_ net48 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1308 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1309 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1310 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1311 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1312 net112 clknet_1_0__leaf__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1313 VGND clknet_1_0__leaf__0462_ net112 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1314 net112 clknet_1_0__leaf__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1315 VPWR clknet_1_0__leaf__0462_ net112 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1316 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1317 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1318 net126 clknet_1_0__leaf__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1319 VGND clknet_1_0__leaf__0463_ net126 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1320 net126 clknet_1_0__leaf__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1321 VPWR clknet_1_0__leaf__0463_ net126 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1322 VPWR net35 hold12/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1323 VGND hold12/a_285_47# hold12/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1324 net159 hold12/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1325 VGND net35 hold12/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1326 VPWR hold12/a_285_47# hold12/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1327 hold12/a_285_47# hold12/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1328 hold12/a_285_47# hold12/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1329 net159 hold12/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1330 VPWR acc0.A\[3\] hold23/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1331 VGND hold23/a_285_47# hold23/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1332 net170 hold23/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1333 VGND acc0.A\[3\] hold23/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1334 VPWR hold23/a_285_47# hold23/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1335 hold23/a_285_47# hold23/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1336 hold23/a_285_47# hold23/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1337 net170 hold23/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1338 VPWR acc0.A\[9\] hold34/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1339 VGND hold34/a_285_47# hold34/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1340 net181 hold34/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1341 VGND acc0.A\[9\] hold34/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1342 VPWR hold34/a_285_47# hold34/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1343 hold34/a_285_47# hold34/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1344 hold34/a_285_47# hold34/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1345 net181 hold34/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1346 VPWR acc0.A\[11\] hold45/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1347 VGND hold45/a_285_47# hold45/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1348 net192 hold45/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1349 VGND acc0.A\[11\] hold45/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1350 VPWR hold45/a_285_47# hold45/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1351 hold45/a_285_47# hold45/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1352 hold45/a_285_47# hold45/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1353 net192 hold45/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1354 VPWR comp0.B\[2\] hold56/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1355 VGND hold56/a_285_47# hold56/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1356 net203 hold56/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1357 VGND comp0.B\[2\] hold56/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1358 VPWR hold56/a_285_47# hold56/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1359 hold56/a_285_47# hold56/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1360 hold56/a_285_47# hold56/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1361 net203 hold56/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1362 VPWR net66 hold67/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1363 VGND hold67/a_285_47# hold67/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1364 net214 hold67/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1365 VGND net66 hold67/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1366 VPWR hold67/a_285_47# hold67/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1367 hold67/a_285_47# hold67/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1368 hold67/a_285_47# hold67/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1369 net214 hold67/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1370 VPWR net60 hold78/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1371 VGND hold78/a_285_47# hold78/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1372 net225 hold78/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1373 VGND net60 hold78/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1374 VPWR hold78/a_285_47# hold78/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1375 hold78/a_285_47# hold78/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1376 hold78/a_285_47# hold78/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1377 net225 hold78/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1378 VPWR control0.state\[2\] hold89/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1379 VGND hold89/a_285_47# hold89/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1380 net236 hold89/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1381 VGND control0.state\[2\] hold89/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1382 VPWR hold89/a_285_47# hold89/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1383 hold89/a_285_47# hold89/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1384 hold89/a_285_47# hold89/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1385 net236 hold89/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1386 net45 _1000_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1387 _1000_/a_891_413# _1000_/a_193_47# _1000_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X1388 _1000_/a_561_413# _1000_/a_27_47# _1000_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X1389 VPWR net86 _1000_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1390 net45 _1000_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1391 _1000_/a_381_47# _0098_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X1392 VGND _1000_/a_634_159# _1000_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X1393 VPWR _1000_/a_891_413# _1000_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1394 _1000_/a_466_413# _1000_/a_193_47# _1000_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1395 VPWR _1000_/a_634_159# _1000_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1396 _1000_/a_634_159# _1000_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X1397 _1000_/a_634_159# _1000_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X1398 _1000_/a_975_413# _1000_/a_193_47# _1000_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X1399 VGND _1000_/a_1059_315# _1000_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X1400 _1000_/a_193_47# _1000_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X1401 _1000_/a_891_413# _1000_/a_27_47# _1000_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1402 _1000_/a_592_47# _1000_/a_193_47# _1000_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X1403 VPWR _1000_/a_1059_315# _1000_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1404 _1000_/a_1017_47# _1000_/a_27_47# _1000_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X1405 _1000_/a_193_47# _1000_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X1406 _1000_/a_466_413# _1000_/a_27_47# _1000_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X1407 VGND _1000_/a_891_413# _1000_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1408 _1000_/a_381_47# _0098_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1409 VGND net86 _1000_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1410 VPWR _0343_ _0715_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X1411 VGND _0715_/a_27_47# _0346_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X1412 VGND _0715_/a_27_47# _0346_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1413 _0346_ _0715_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X1414 _0346_ _0715_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1415 VGND _0343_ _0715_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X1416 VPWR _0715_/a_27_47# _0346_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1417 _0346_ _0715_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1418 _0346_ _0715_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1419 VPWR _0715_/a_27_47# _0346_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1420 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X1421 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X1422 VPWR _0183_ _0577_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X1423 _0577_/a_27_297# _0217_ _0577_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X1424 VGND _0183_ _0577_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X1425 _0120_ _0577_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1426 _0577_/a_27_297# _0217_ _0577_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X1427 _0577_/a_109_297# acc0.A\[22\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1428 _0577_/a_373_47# acc0.A\[22\] _0577_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1429 _0120_ _0577_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1430 _0577_/a_109_297# net150 _0577_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1431 _0577_/a_109_47# net150 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1432 _0646_/a_377_297# acc0.A\[13\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=2.42 as=0 ps=0 w=1 l=0.15
X1433 _0646_/a_47_47# net40 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1434 _0646_/a_129_47# net40 _0646_/a_47_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.72 as=0.169 ps=1.82 w=0.65 l=0.15
X1435 _0646_/a_285_47# net40 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X1436 _0278_ _0646_/a_47_47# _0646_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X1437 VGND acc0.A\[13\] _0646_/a_129_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1438 VPWR acc0.A\[13\] _0646_/a_47_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1439 VPWR _0646_/a_47_47# _0278_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.33 ps=2.66 w=1 l=0.15
X1440 _0278_ net40 _0646_/a_377_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1441 _0646_/a_285_47# acc0.A\[13\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1442 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X1443 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X1444 VPWR output57/a_27_47# pp[29] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1445 pp[29] output57/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1446 VPWR net57 output57/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1447 pp[29] output57/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X1448 VGND output57/a_27_47# pp[29] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1449 VGND net57 output57/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1450 VPWR output46/a_27_47# pp[19] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1451 pp[19] output46/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1452 VPWR net46 output46/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1453 pp[19] output46/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X1454 VGND output46/a_27_47# pp[19] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1455 VGND net46 output46/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1456 VPWR output35/a_27_47# done VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1457 done output35/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1458 VPWR net35 output35/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1459 done output35/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X1460 VGND output35/a_27_47# done VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1461 VGND net35 output35/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1462 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1463 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1464 VPWR _0178_ _0500_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X1465 VGND _0500_/a_27_47# _0179_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X1466 VGND _0500_/a_27_47# _0179_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1467 _0179_ _0500_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X1468 _0179_ _0500_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1469 VGND _0178_ _0500_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X1470 VPWR _0500_/a_27_47# _0179_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1471 _0179_ _0500_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1472 _0179_ _0500_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1473 VPWR _0500_/a_27_47# _0179_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1474 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1475 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1476 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1477 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1478 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1479 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1480 VPWR net58 _0629_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X1481 _0261_ _0629_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X1482 VGND net58 _0629_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X1483 _0629_/a_59_75# acc0.A\[2\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1484 _0261_ _0629_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X1485 _0629_/a_145_75# acc0.A\[2\] _0629_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X1486 _0490_ _0483_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1487 VGND _0483_ _0490_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1488 _0490_ _0483_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1489 VPWR _0483_ _0490_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1490 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1491 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1492 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1493 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1494 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1495 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1496 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1497 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1498 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X1499 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X1500 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1501 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1502 _0481_ _0963_/a_35_297# _0963_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1503 _0481_ control0.count\[0\] _0963_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X1504 _0963_/a_35_297# control0.count\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1505 _0963_/a_117_297# control0.count\[0\] _0963_/a_35_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1506 VPWR control0.count\[0\] _0963_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1507 VGND control0.count\[1\] _0963_/a_35_297# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1508 VGND _0963_/a_35_297# _0481_ VGND sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X1509 _0963_/a_285_297# control0.count\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1510 VPWR control0.count\[1\] _0963_/a_117_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1511 _0963_/a_285_47# control0.count\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1512 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1513 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1514 VPWR _0946_/a_30_53# _0466_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.315 pd=2.63 as=0.135 ps=1.27 w=1 l=0.15
X1515 VGND _0946_/a_30_53# _0466_ VGND sky130_fd_pr__nfet_01v8 ad=0.18525 pd=1.87 as=0.08775 ps=0.92 w=0.65 l=0.15
X1516 _0466_ _0946_/a_30_53# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14825 ps=1.34 w=1 l=0.15
X1517 _0946_/a_112_297# control0.state\[0\] _0946_/a_30_53# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1518 _0466_ _0946_/a_30_53# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10187 ps=0.99 w=0.65 l=0.15
X1519 VGND net34 _0946_/a_30_53# VGND sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1520 _0946_/a_30_53# control0.state\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1521 VGND control0.state\[0\] _0946_/a_30_53# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1522 _0946_/a_184_297# control0.state\[1\] _0946_/a_112_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1523 VPWR net34 _0946_/a_184_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1524 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X1525 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X1526 clkload1/Y clknet_1_0__leaf__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.25
X1527 VGND clknet_1_0__leaf__0465_ clkload1/a_268_47# VGND sky130_fd_pr__nfet_01v8 ad=0.14575 pd=1.63 as=0.05775 ps=0.76 w=0.55 l=0.15
X1528 clkload1/Y clknet_1_0__leaf__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X1529 clkload1/Y clknet_1_0__leaf__0465_ clkload1/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0.077 pd=0.83 as=0.05775 ps=0.76 w=0.55 l=0.15
X1530 VPWR clknet_1_0__leaf__0465_ clkload1/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.25
X1531 clkload1/a_110_47# clknet_1_0__leaf__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.76 as=0.14575 ps=1.63 w=0.55 l=0.15
X1532 clkload1/a_268_47# clknet_1_0__leaf__0465_ clkload1/Y VGND sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.76 as=0.077 ps=0.83 w=0.55 l=0.15
X1533 VPWR clknet_1_0__leaf__0465_ clkload1/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.25
X1534 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1535 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1536 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1537 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1538 _0800_/a_240_47# net245 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1539 _0093_ _0800_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1540 VGND _0219_ _0800_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1541 _0800_/a_51_297# _0413_ _0800_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.4125 pd=1.825 as=0.105 ps=1.21 w=1 l=0.15
X1542 _0800_/a_149_47# _0345_ _0800_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.09912 pd=0.955 as=0.2015 ps=1.92 w=0.65 l=0.15
X1543 _0800_/a_240_47# _0412_ _0800_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.09912 ps=0.955 w=0.65 l=0.15
X1544 VPWR _0219_ _0800_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.105 ps=1.21 w=1 l=0.15
X1545 _0093_ _0800_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.165 ps=1.33 w=1 l=0.15
X1546 _0800_/a_149_47# _0413_ _0800_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1547 _0800_/a_245_297# _0412_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X1548 VPWR _0345_ _0800_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.34 ps=2.68 w=1 l=0.15
X1549 _0800_/a_512_297# net245 _0800_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.4125 ps=1.825 w=1 l=0.15
X1550 _0731_/a_81_21# _0326_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X1551 _0731_/a_299_297# _0326_ _0731_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X1552 VPWR _0731_/a_81_21# _0359_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1553 VPWR _0250_ _0731_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1554 VGND _0731_/a_81_21# _0359_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1555 VGND _0312_ _0731_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X1556 _0731_/a_299_297# _0312_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1557 _0731_/a_384_47# _0250_ _0731_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1558 VPWR _0222_ _0225_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1559 _0225_ _0222_ _0593_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X1560 _0593_/a_113_47# _0224_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1561 _0225_ _0224_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1562 _0662_/a_81_21# _0293_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X1563 _0662_/a_299_297# _0293_ _0662_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X1564 VPWR _0662_/a_81_21# _0294_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1565 VPWR _0259_ _0662_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1566 VGND _0662_/a_81_21# _0294_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1567 VGND _0275_ _0662_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X1568 _0662_/a_299_297# _0275_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1569 _0662_/a_384_47# _0259_ _0662_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1570 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1571 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1572 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1573 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1574 VPWR comp0.B\[5\] hold13/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1575 VGND hold13/a_285_47# hold13/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1576 net160 hold13/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1577 VGND comp0.B\[5\] hold13/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1578 VPWR hold13/a_285_47# hold13/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1579 hold13/a_285_47# hold13/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1580 hold13/a_285_47# hold13/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1581 net160 hold13/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1582 VPWR comp0.B\[7\] hold24/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1583 VGND hold24/a_285_47# hold24/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1584 net171 hold24/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1585 VGND comp0.B\[7\] hold24/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1586 VPWR hold24/a_285_47# hold24/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1587 hold24/a_285_47# hold24/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1588 hold24/a_285_47# hold24/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1589 net171 hold24/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1590 VPWR _0154_ hold35/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1591 VGND hold35/a_285_47# hold35/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1592 net182 hold35/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1593 VGND _0154_ hold35/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1594 VPWR hold35/a_285_47# hold35/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1595 hold35/a_285_47# hold35/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1596 hold35/a_285_47# hold35/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1597 net182 hold35/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1598 VPWR comp0.B\[13\] hold46/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1599 VGND hold46/a_285_47# hold46/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1600 net193 hold46/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1601 VGND comp0.B\[13\] hold46/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1602 VPWR hold46/a_285_47# hold46/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1603 hold46/a_285_47# hold46/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1604 hold46/a_285_47# hold46/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1605 net193 hold46/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1606 VPWR comp0.B\[6\] hold57/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1607 VGND hold57/a_285_47# hold57/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1608 net204 hold57/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1609 VGND comp0.B\[6\] hold57/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1610 VPWR hold57/a_285_47# hold57/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1611 hold57/a_285_47# hold57/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1612 hold57/a_285_47# hold57/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1613 net204 hold57/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1614 VPWR acc0.A\[23\] hold68/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1615 VGND hold68/a_285_47# hold68/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1616 net215 hold68/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1617 VGND acc0.A\[23\] hold68/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1618 VPWR hold68/a_285_47# hold68/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1619 hold68/a_285_47# hold68/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1620 hold68/a_285_47# hold68/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1621 net215 hold68/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1622 VPWR control0.count\[1\] hold79/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1623 VGND hold79/a_285_47# hold79/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1624 net226 hold79/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1625 VGND control0.count\[1\] hold79/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1626 VPWR hold79/a_285_47# hold79/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1627 hold79/a_285_47# hold79/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1628 hold79/a_285_47# hold79/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1629 net226 hold79/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1630 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X1631 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X1632 _0714_/a_240_47# _0219_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X1633 _0111_ _0714_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X1634 VGND net225 _0714_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1635 _0714_/a_51_297# _0344_ _0714_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X1636 _0714_/a_149_47# _0345_ _0714_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X1637 _0714_/a_240_47# _0342_ _0714_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1638 VPWR net225 _0714_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X1639 _0111_ _0714_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X1640 _0714_/a_149_47# _0344_ _0714_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1641 _0714_/a_245_297# _0342_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1642 VPWR _0345_ _0714_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1643 _0714_/a_512_297# _0219_ _0714_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1644 _0645_/a_377_297# acc0.A\[14\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=2.42 as=0 ps=0 w=1 l=0.15
X1645 _0645_/a_47_47# net41 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1646 _0645_/a_129_47# net41 _0645_/a_47_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.72 as=0.169 ps=1.82 w=0.65 l=0.15
X1647 _0645_/a_285_47# net41 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X1648 _0277_ _0645_/a_47_47# _0645_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X1649 VGND acc0.A\[14\] _0645_/a_129_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1650 VPWR acc0.A\[14\] _0645_/a_47_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1651 VPWR _0645_/a_47_47# _0277_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.33 ps=2.66 w=1 l=0.15
X1652 _0277_ net41 _0645_/a_377_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1653 _0645_/a_285_47# acc0.A\[14\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1654 VPWR _0183_ _0576_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X1655 _0576_/a_27_297# _0217_ _0576_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X1656 VGND _0183_ _0576_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X1657 _0121_ _0576_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1658 _0576_/a_27_297# _0217_ _0576_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X1659 _0576_/a_109_297# acc0.A\[23\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1660 _0576_/a_373_47# acc0.A\[23\] _0576_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1661 _0121_ _0576_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1662 _0576_/a_109_297# net176 _0576_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1663 _0576_/a_109_47# net176 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1664 acc0.A\[13\] _1059_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1665 _1059_/a_891_413# _1059_/a_193_47# _1059_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X1666 _1059_/a_561_413# _1059_/a_27_47# _1059_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X1667 VPWR net145 _1059_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1668 acc0.A\[13\] _1059_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1669 _1059_/a_381_47# _0157_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X1670 VGND _1059_/a_634_159# _1059_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X1671 VPWR _1059_/a_891_413# _1059_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1672 _1059_/a_466_413# _1059_/a_193_47# _1059_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1673 VPWR _1059_/a_634_159# _1059_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1674 _1059_/a_634_159# _1059_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X1675 _1059_/a_634_159# _1059_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X1676 _1059_/a_975_413# _1059_/a_193_47# _1059_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X1677 VGND _1059_/a_1059_315# _1059_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X1678 _1059_/a_193_47# _1059_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X1679 _1059_/a_891_413# _1059_/a_27_47# _1059_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1680 _1059_/a_592_47# _1059_/a_193_47# _1059_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X1681 VPWR _1059_/a_1059_315# _1059_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1682 _1059_/a_1017_47# _1059_/a_27_47# _1059_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X1683 _1059_/a_193_47# _1059_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X1684 _1059_/a_466_413# _1059_/a_27_47# _1059_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X1685 VGND _1059_/a_891_413# _1059_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1686 _1059_/a_381_47# _0157_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1687 VGND net145 _1059_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1688 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X1689 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X1690 VPWR output36/a_27_47# pp[0] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1691 pp[0] output36/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1692 VPWR net36 output36/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1693 pp[0] output36/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X1694 VGND output36/a_27_47# pp[0] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1695 VGND net36 output36/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1696 VPWR net58 output58/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X1697 VGND output58/a_27_47# pp[2] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X1698 VGND output58/a_27_47# pp[2] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1699 pp[2] output58/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X1700 pp[2] output58/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1701 VGND net58 output58/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X1702 VPWR output58/a_27_47# pp[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1703 pp[2] output58/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1704 pp[2] output58/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1705 VPWR output58/a_27_47# pp[2] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1706 VPWR net47 output47/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X1707 VGND output47/a_27_47# pp[1] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X1708 VGND output47/a_27_47# pp[1] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1709 pp[1] output47/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X1710 pp[1] output47/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1711 VGND net47 output47/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X1712 VPWR output47/a_27_47# pp[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1713 pp[1] output47/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1714 pp[1] output47/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1715 VPWR output47/a_27_47# pp[1] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1716 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1717 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1718 net104 clknet_1_0__leaf__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1719 VGND clknet_1_0__leaf__0461_ net104 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1720 net104 clknet_1_0__leaf__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1721 VPWR clknet_1_0__leaf__0461_ net104 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1722 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1723 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1724 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1725 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1726 VPWR acc0.A\[3\] _0628_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X1727 VGND acc0.A\[3\] _0260_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1728 _0628_/a_109_297# net61 _0260_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1729 _0260_ net61 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1730 _0559_/a_240_47# net26 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X1731 _0133_ _0559_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X1732 VGND _0208_ _0559_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1733 _0559_/a_51_297# net205 _0559_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X1734 _0559_/a_149_47# _0212_ _0559_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X1735 _0559_/a_240_47# _0173_ _0559_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1736 VPWR _0208_ _0559_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X1737 _0133_ _0559_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X1738 _0559_/a_149_47# net205 _0559_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1739 _0559_/a_245_297# _0173_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1740 VPWR _0212_ _0559_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1741 _0559_/a_512_297# net26 _0559_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1742 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1743 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1744 net85 clknet_1_1__leaf__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1745 VGND clknet_1_1__leaf__0459_ net85 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1746 net85 clknet_1_1__leaf__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1747 VPWR clknet_1_1__leaf__0459_ net85 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1748 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1749 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1750 VPWR _0478_ _0962_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X1751 VGND _0478_ _0480_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1752 _0962_/a_109_297# _0479_ _0480_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1753 _0480_ _0479_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1754 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1755 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1756 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1757 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1758 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X1759 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X1760 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X1761 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X1762 clkload2/Y clknet_1_0__leaf__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.25
X1763 VGND clknet_1_0__leaf__0464_ clkload2/a_268_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1155 ps=1.52 w=0.55 l=0.15
X1764 clkload2/Y clknet_1_0__leaf__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.25
X1765 clkload2/Y clknet_1_0__leaf__0464_ clkload2/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0.154 pd=1.66 as=0.1155 ps=1.52 w=0.55 l=0.15
X1766 VPWR clknet_1_0__leaf__0464_ clkload2/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.25
X1767 clkload2/a_110_47# clknet_1_0__leaf__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.15
X1768 clkload2/a_268_47# clknet_1_0__leaf__0464_ clkload2/Y VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.15
X1769 VPWR clknet_1_0__leaf__0464_ clkload2/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.25
X1770 _0661_/a_27_297# _0288_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.252 pd=2.88 as=0 ps=0 w=0.42 l=0.15
X1771 _0661_/a_27_297# _0292_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1772 _0661_/a_277_297# _0288_ _0661_/a_205_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1386 pd=1.5 as=0.0882 ps=1.26 w=0.42 l=0.15
X1773 VPWR _0287_ _0661_/a_277_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1774 _0293_ _0661_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X1775 _0661_/a_205_297# _0289_ _0661_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1386 ps=1.5 w=0.42 l=0.15
X1776 _0293_ _0661_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1777 VGND _0289_ _0661_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1778 _0661_/a_109_297# _0292_ _0661_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1779 VGND _0287_ _0661_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1780 VGND _0347_ _0730_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X1781 _0730_/a_510_47# _0358_ _0730_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X1782 _0730_/a_79_21# _0352_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X1783 VPWR _0358_ _0730_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1784 _0730_/a_79_21# _0357_ _0730_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X1785 _0730_/a_297_297# _0347_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1786 _0730_/a_79_21# _0352_ _0730_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X1787 VPWR _0730_/a_79_21# _0108_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1788 VGND _0730_/a_79_21# _0108_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1789 _0730_/a_215_47# _0357_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1790 VGND acc0.A\[22\] _0592_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X1791 _0592_/a_68_297# net50 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1792 _0224_ _0592_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1793 VPWR acc0.A\[22\] _0592_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X1794 _0224_ _0592_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X1795 _0592_/a_150_297# net50 _0592_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1796 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X1797 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X1798 VPWR _0134_ hold14/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1799 VGND hold14/a_285_47# hold14/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1800 net161 hold14/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1801 VGND _0134_ hold14/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1802 VPWR hold14/a_285_47# hold14/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1803 hold14/a_285_47# hold14/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1804 hold14/a_285_47# hold14/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1805 net161 hold14/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1806 VPWR _0136_ hold25/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1807 VGND hold25/a_285_47# hold25/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1808 net172 hold25/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1809 VGND _0136_ hold25/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1810 VPWR hold25/a_285_47# hold25/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1811 hold25/a_285_47# hold25/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1812 hold25/a_285_47# hold25/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1813 net172 hold25/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1814 VPWR comp0.B\[14\] hold36/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1815 VGND hold36/a_285_47# hold36/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1816 net183 hold36/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1817 VGND comp0.B\[14\] hold36/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1818 VPWR hold36/a_285_47# hold36/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1819 hold36/a_285_47# hold36/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1820 hold36/a_285_47# hold36/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1821 net183 hold36/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1822 VPWR _0142_ hold47/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1823 VGND hold47/a_285_47# hold47/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1824 net194 hold47/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1825 VGND _0142_ hold47/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1826 VPWR hold47/a_285_47# hold47/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1827 hold47/a_285_47# hold47/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1828 hold47/a_285_47# hold47/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1829 net194 hold47/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1830 VPWR comp0.B\[4\] hold58/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1831 VGND hold58/a_285_47# hold58/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1832 net205 hold58/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1833 VGND comp0.B\[4\] hold58/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1834 VPWR hold58/a_285_47# hold58/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1835 hold58/a_285_47# hold58/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1836 hold58/a_285_47# hold58/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1837 net205 hold58/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1838 VPWR net52 hold69/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1839 VGND hold69/a_285_47# hold69/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1840 net216 hold69/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1841 VGND net52 hold69/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1842 VPWR hold69/a_285_47# hold69/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1843 hold69/a_285_47# hold69/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1844 hold69/a_285_47# hold69/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1845 net216 hold69/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1846 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1847 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1848 net117 clknet_1_1__leaf__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1849 VGND clknet_1_1__leaf__0462_ net117 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1850 net117 clknet_1_1__leaf__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1851 VPWR clknet_1_1__leaf__0462_ net117 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1852 VPWR _0208_ _0713_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X1853 VGND _0713_/a_27_47# _0345_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X1854 VGND _0713_/a_27_47# _0345_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1855 _0345_ _0713_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X1856 _0345_ _0713_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1857 VGND _0208_ _0713_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X1858 VPWR _0713_/a_27_47# _0345_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1859 _0345_ _0713_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1860 _0345_ _0713_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1861 VPWR _0713_/a_27_47# _0345_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1862 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1863 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1864 _0644_/a_377_297# acc0.A\[15\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=2.42 as=0 ps=0 w=1 l=0.15
X1865 _0644_/a_47_47# net42 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1866 _0644_/a_129_47# net42 _0644_/a_47_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.72 as=0.169 ps=1.82 w=0.65 l=0.15
X1867 _0644_/a_285_47# net42 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X1868 _0276_ _0644_/a_47_47# _0644_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X1869 VGND acc0.A\[15\] _0644_/a_129_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1870 VPWR acc0.A\[15\] _0644_/a_47_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1871 VPWR _0644_/a_47_47# _0276_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.33 ps=2.66 w=1 l=0.15
X1872 _0276_ net42 _0644_/a_377_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1873 _0644_/a_285_47# acc0.A\[15\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1874 VPWR _0216_ _0575_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X1875 _0575_/a_27_297# _0217_ _0575_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X1876 VGND _0216_ _0575_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X1877 _0122_ _0575_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1878 _0575_/a_27_297# _0217_ _0575_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X1879 _0575_/a_109_297# net199 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1880 _0575_/a_373_47# net199 _0575_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1881 _0122_ _0575_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1882 _0575_/a_109_297# net215 _0575_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1883 _0575_/a_109_47# net215 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1884 acc0.A\[12\] _1058_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1885 _1058_/a_891_413# _1058_/a_193_47# _1058_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X1886 _1058_/a_561_413# _1058_/a_27_47# _1058_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X1887 VPWR net144 _1058_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1888 acc0.A\[12\] _1058_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1889 _1058_/a_381_47# _0156_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X1890 VGND _1058_/a_634_159# _1058_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X1891 VPWR _1058_/a_891_413# _1058_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1892 _1058_/a_466_413# _1058_/a_193_47# _1058_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1893 VPWR _1058_/a_634_159# _1058_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1894 _1058_/a_634_159# _1058_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X1895 _1058_/a_634_159# _1058_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X1896 _1058_/a_975_413# _1058_/a_193_47# _1058_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X1897 VGND _1058_/a_1059_315# _1058_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X1898 _1058_/a_193_47# _1058_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X1899 _1058_/a_891_413# _1058_/a_27_47# _1058_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1900 _1058_/a_592_47# _1058_/a_193_47# _1058_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X1901 VPWR _1058_/a_1059_315# _1058_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1902 _1058_/a_1017_47# _1058_/a_27_47# _1058_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X1903 _1058_/a_193_47# _1058_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X1904 _1058_/a_466_413# _1058_/a_27_47# _1058_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X1905 VGND _1058_/a_891_413# _1058_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X1906 _1058_/a_381_47# _0156_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1907 VGND net144 _1058_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1908 VPWR output59/a_27_47# pp[30] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1909 pp[30] output59/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1910 VPWR net59 output59/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1911 pp[30] output59/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X1912 VGND output59/a_27_47# pp[30] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1913 VGND net59 output59/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1914 VPWR output48/a_27_47# pp[20] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1915 pp[20] output48/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1916 VPWR net48 output48/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X1917 pp[20] output48/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X1918 VGND output48/a_27_47# pp[20] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1919 VGND net48 output48/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1920 VPWR net37 output37/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X1921 VGND output37/a_27_47# pp[10] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X1922 VGND output37/a_27_47# pp[10] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1923 pp[10] output37/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X1924 pp[10] output37/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1925 VGND net37 output37/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X1926 VPWR output37/a_27_47# pp[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1927 pp[10] output37/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1928 pp[10] output37/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1929 VPWR output37/a_27_47# pp[10] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1930 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1931 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1932 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X1933 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X1934 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1935 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1936 _0627_/a_109_93# _0258_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1937 _0627_/a_215_53# _0255_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1938 VGND _0627_/a_109_93# _0627_/a_215_53# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1939 VGND _0254_ _0627_/a_215_53# VGND sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1940 VPWR _0254_ _0627_/a_369_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06825 ps=0.745 w=0.42 l=0.15
X1941 _0627_/a_369_297# _0255_ _0627_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.0441 ps=0.63 w=0.42 l=0.15
X1942 _0259_ _0627_/a_215_53# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X1943 _0627_/a_297_297# _0627_/a_109_93# _0627_/a_215_53# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1944 _0627_/a_109_93# _0258_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1945 _0259_ _0627_/a_215_53# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10025 ps=0.985 w=0.65 l=0.15
X1946 VGND net185 _0558_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X1947 _0558_/a_68_297# _0175_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X1948 _0212_ _0558_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1949 VPWR net185 _0558_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X1950 _0212_ _0558_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X1951 _0558_/a_150_297# _0175_ _0558_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1952 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1953 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1954 VPWR acc0.A\[14\] hold100/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1955 VGND hold100/a_285_47# hold100/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1956 net247 hold100/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X1957 VGND acc0.A\[14\] hold100/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X1958 VPWR hold100/a_285_47# hold100/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X1959 hold100/a_285_47# hold100/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1960 hold100/a_285_47# hold100/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X1961 net247 hold100/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X1962 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X1963 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X1964 net89 clknet_1_0__leaf__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1965 VGND clknet_1_0__leaf__0460_ net89 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1966 net89 clknet_1_0__leaf__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1967 VPWR clknet_1_0__leaf__0460_ net89 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1968 _0961_/a_199_47# control0.count\[1\] _0479_ VGND sky130_fd_pr__nfet_01v8 ad=0.09588 pd=0.945 as=0.091 ps=0.93 w=0.65 l=0.15
X1969 _0961_/a_113_297# control0.count\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.1475 ps=1.295 w=1 l=0.15
X1970 _0479_ control0.count\[2\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.17225 ps=1.83 w=0.65 l=0.15
X1971 VPWR control0.count\[1\] _0961_/a_113_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1475 pd=1.295 as=0.14 ps=1.28 w=1 l=0.15
X1972 _0961_/a_113_297# control0.count\[2\] _0479_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X1973 VGND control0.count\[0\] _0961_/a_199_47# VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.09588 ps=0.945 w=0.65 l=0.15
X1974 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X1975 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X1976 net123 clknet_1_0__leaf__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X1977 VGND clknet_1_0__leaf__0463_ net123 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1978 net123 clknet_1_0__leaf__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1979 VPWR clknet_1_0__leaf__0463_ net123 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1980 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X1981 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X1982 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X1983 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X1984 clkload3/Y clknet_1_1__leaf__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.25
X1985 VGND clknet_1_1__leaf__0461_ clkload3/a_268_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1155 ps=1.52 w=0.55 l=0.15
X1986 clkload3/Y clknet_1_1__leaf__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.25
X1987 clkload3/Y clknet_1_1__leaf__0461_ clkload3/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0.154 pd=1.66 as=0.1155 ps=1.52 w=0.55 l=0.15
X1988 VPWR clknet_1_1__leaf__0461_ clkload3/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.25
X1989 clkload3/a_110_47# clknet_1_1__leaf__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.15
X1990 clkload3/a_268_47# clknet_1_1__leaf__0461_ clkload3/Y VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.15
X1991 VPWR clknet_1_1__leaf__0461_ clkload3/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.25
X1992 VPWR _0290_ _0292_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X1993 _0292_ _0290_ _0660_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X1994 _0660_/a_113_47# _0291_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X1995 _0292_ _0291_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X1996 VPWR acc0.A\[23\] _0591_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X1997 VGND acc0.A\[23\] _0223_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X1998 _0591_/a_109_297# net51 _0223_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X1999 _0223_ net51 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2000 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2001 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2002 _0789_/a_75_199# _0277_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13487 ps=1.065 w=0.65 l=0.15
X2003 _0789_/a_208_47# _0404_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.12513 pd=1.035 as=0.11213 ps=0.995 w=0.65 l=0.15
X2004 _0789_/a_315_47# _0298_ _0789_/a_208_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.17 as=0.12513 ps=1.035 w=0.65 l=0.15
X2005 VGND _0297_ _0789_/a_75_199# VGND sky130_fd_pr__nfet_01v8 ad=0.13487 pd=1.065 as=0.10563 ps=0.975 w=0.65 l=0.15
X2006 _0789_/a_75_199# _0299_ _0789_/a_315_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10563 pd=0.975 as=0.169 ps=1.17 w=0.65 l=0.15
X2007 _0789_/a_75_199# _0277_ _0789_/a_544_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2075 ps=1.415 w=1 l=0.15
X2008 _0789_/a_544_297# _0297_ _0789_/a_201_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2075 pd=1.415 as=0.1625 ps=1.325 w=1 l=0.15
X2009 VPWR _0789_/a_75_199# _0405_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1425 pd=1.285 as=0.285 ps=2.57 w=1 l=0.15
X2010 _0789_/a_201_297# _0404_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.1425 ps=1.285 w=1 l=0.15
X2011 VPWR _0298_ _0789_/a_201_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.305 pd=1.61 as=0.165 ps=1.33 w=1 l=0.15
X2012 _0789_/a_201_297# _0299_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.305 ps=1.61 w=1 l=0.15
X2013 VGND _0789_/a_75_199# _0405_ VGND sky130_fd_pr__nfet_01v8 ad=0.11213 pd=0.995 as=0.169 ps=1.82 w=0.65 l=0.15
X2014 VPWR clknet_1_1__leaf__0457_ _0858_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2015 _0458_ _0858_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2016 _0458_ _0858_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2017 VGND clknet_1_1__leaf__0457_ _0858_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2018 VPWR acc0.A\[31\] hold15/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2019 VGND hold15/a_285_47# hold15/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2020 net162 hold15/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2021 VGND acc0.A\[31\] hold15/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2022 VPWR hold15/a_285_47# hold15/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2023 hold15/a_285_47# hold15/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2024 hold15/a_285_47# hold15/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2025 net162 hold15/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2026 VPWR comp0.B\[9\] hold26/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2027 VGND hold26/a_285_47# hold26/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2028 net173 hold26/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2029 VGND comp0.B\[9\] hold26/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2030 VPWR hold26/a_285_47# hold26/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2031 hold26/a_285_47# hold26/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2032 hold26/a_285_47# hold26/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2033 net173 hold26/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2034 VPWR _0143_ hold37/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2035 VGND hold37/a_285_47# hold37/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2036 net184 hold37/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2037 VGND _0143_ hold37/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2038 VPWR hold37/a_285_47# hold37/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2039 hold37/a_285_47# hold37/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2040 hold37/a_285_47# hold37/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2041 net184 hold37/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2042 VPWR comp0.B\[12\] hold48/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2043 VGND hold48/a_285_47# hold48/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2044 net195 hold48/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2045 VGND comp0.B\[12\] hold48/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2046 VPWR hold48/a_285_47# hold48/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2047 hold48/a_285_47# hold48/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2048 hold48/a_285_47# hold48/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2049 net195 hold48/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2050 VPWR acc0.A\[18\] hold59/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2051 VGND hold59/a_285_47# hold59/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2052 net206 hold59/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2053 VGND acc0.A\[18\] hold59/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2054 VPWR hold59/a_285_47# hold59/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2055 hold59/a_285_47# hold59/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2056 hold59/a_285_47# hold59/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2057 net206 hold59/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2058 net73 clknet_1_1__leaf__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2059 VGND clknet_1_1__leaf__0458_ net73 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2060 net73 clknet_1_1__leaf__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2061 VPWR clknet_1_1__leaf__0458_ net73 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2062 _0643_/a_103_199# _0274_ _0643_/a_253_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X2063 VPWR _0643_/a_103_199# _0275_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X2064 _0643_/a_337_297# _0269_ _0643_/a_253_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2065 _0643_/a_103_199# _0272_ _0643_/a_337_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.165 ps=1.33 w=1 l=0.15
X2066 _0643_/a_253_297# _0260_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X2067 VPWR _0274_ _0643_/a_103_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.2125 ps=1.425 w=1 l=0.15
X2068 VGND _0643_/a_103_199# _0275_ VGND sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X2069 _0643_/a_253_47# _0260_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12675 ps=1.04 w=0.65 l=0.15
X2070 _0643_/a_253_47# _0272_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X2071 VGND _0269_ _0643_/a_253_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X2072 _0712_/a_465_47# _0339_ _0712_/a_381_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.1755 ps=1.84 w=0.65 l=0.15
X2073 VGND _0341_ _0712_/a_561_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2145 ps=1.96 w=0.65 l=0.15
X2074 VPWR _0340_ _0712_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.86 ps=7.72 w=1 l=0.15
X2075 _0712_/a_297_297# _0339_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2076 _0712_/a_297_297# _0341_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2077 VPWR _0220_ _0712_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2078 _0712_/a_381_47# _0220_ _0712_/a_79_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.36725 ps=2.43 w=0.65 l=0.15
X2079 _0712_/a_297_297# _0343_ _0712_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2080 VPWR _0712_/a_79_21# _0344_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2081 _0712_/a_79_21# _0343_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2082 VGND _0712_/a_79_21# _0344_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2083 _0712_/a_561_47# _0340_ _0712_/a_465_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2084 VPWR _0216_ _0574_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X2085 _0574_/a_27_297# _0217_ _0574_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X2086 VGND _0216_ _0574_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X2087 _0123_ _0574_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2088 _0574_/a_27_297# _0217_ _0574_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X2089 _0574_/a_109_297# acc0.A\[25\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2090 _0574_/a_373_47# acc0.A\[25\] _0574_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2091 _0123_ _0574_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2092 _0574_/a_109_297# net199 _0574_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2093 _0574_/a_109_47# net199 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2094 acc0.A\[11\] _1057_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2095 _1057_/a_891_413# _1057_/a_193_47# _1057_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2096 _1057_/a_561_413# _1057_/a_27_47# _1057_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2097 VPWR net143 _1057_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2098 acc0.A\[11\] _1057_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2099 _1057_/a_381_47# net189 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2100 VGND _1057_/a_634_159# _1057_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2101 VPWR _1057_/a_891_413# _1057_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2102 _1057_/a_466_413# _1057_/a_193_47# _1057_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2103 VPWR _1057_/a_634_159# _1057_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2104 _1057_/a_634_159# _1057_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2105 _1057_/a_634_159# _1057_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2106 _1057_/a_975_413# _1057_/a_193_47# _1057_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2107 VGND _1057_/a_1059_315# _1057_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2108 _1057_/a_193_47# _1057_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2109 _1057_/a_891_413# _1057_/a_27_47# _1057_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2110 _1057_/a_592_47# _1057_/a_193_47# _1057_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2111 VPWR _1057_/a_1059_315# _1057_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2112 _1057_/a_1017_47# _1057_/a_27_47# _1057_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2113 _1057_/a_193_47# _1057_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2114 _1057_/a_466_413# _1057_/a_27_47# _1057_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2115 VGND _1057_/a_891_413# _1057_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2116 _1057_/a_381_47# net189 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2117 VGND net143 _1057_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2118 VPWR output49/a_27_47# pp[21] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2119 pp[21] output49/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2120 VPWR net49 output49/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2121 pp[21] output49/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X2122 VGND output49/a_27_47# pp[21] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2123 VGND net49 output49/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2124 VPWR output38/a_27_47# pp[11] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2125 pp[11] output38/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2126 VPWR net38 output38/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2127 pp[11] output38/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X2128 VGND output38/a_27_47# pp[11] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2129 VGND net38 output38/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2130 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X2131 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X2132 VPWR clk clkbuf_0_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X2133 VPWR clkbuf_0_clk/a_110_47# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X2134 clknet_0_clk clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2135 clknet_0_clk clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2136 VPWR clkbuf_0_clk/a_110_47# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2137 VPWR clkbuf_0_clk/a_110_47# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2138 clkbuf_0_clk/a_110_47# clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2139 clkbuf_0_clk/a_110_47# clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X2140 VGND clkbuf_0_clk/a_110_47# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X2141 clknet_0_clk clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2142 VGND clkbuf_0_clk/a_110_47# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2143 clkbuf_0_clk/a_110_47# clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2144 VGND clk clkbuf_0_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2145 VGND clkbuf_0_clk/a_110_47# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2146 VPWR clkbuf_0_clk/a_110_47# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2147 clknet_0_clk clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2148 VGND clk clkbuf_0_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2149 VGND clkbuf_0_clk/a_110_47# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2150 VPWR clkbuf_0_clk/a_110_47# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2151 VGND clkbuf_0_clk/a_110_47# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2152 clknet_0_clk clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2153 clkbuf_0_clk/a_110_47# clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2154 VPWR clk clkbuf_0_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2155 VPWR clkbuf_0_clk/a_110_47# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2156 VPWR clkbuf_0_clk/a_110_47# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2157 VGND clkbuf_0_clk/a_110_47# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2158 clknet_0_clk clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2159 VGND clkbuf_0_clk/a_110_47# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2160 VGND clkbuf_0_clk/a_110_47# clknet_0_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2161 clknet_0_clk clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2162 clknet_0_clk clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2163 clknet_0_clk clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2164 clknet_0_clk clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2165 VPWR clkbuf_0_clk/a_110_47# clknet_0_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2166 clknet_0_clk clkbuf_0_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2167 clknet_0_clk clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2168 clknet_0_clk clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2169 clknet_0_clk clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2170 clknet_0_clk clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2171 clknet_0_clk clkbuf_0_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2172 _0557_/a_240_47# net27 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X2173 _0134_ _0557_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X2174 VGND _0208_ _0557_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2175 _0557_/a_51_297# net160 _0557_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X2176 _0557_/a_149_47# _0211_ _0557_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X2177 _0557_/a_240_47# _0173_ _0557_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2178 VPWR _0208_ _0557_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X2179 _0134_ _0557_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X2180 _0557_/a_149_47# net160 _0557_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2181 _0557_/a_245_297# _0173_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2182 VPWR _0211_ _0557_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2183 _0557_/a_512_297# net27 _0557_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2184 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2185 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2186 VGND _0256_ _0626_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2187 _0626_/a_68_297# _0257_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2188 _0258_ _0626_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2189 VPWR _0256_ _0626_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X2190 _0258_ _0626_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X2191 _0626_/a_150_297# _0257_ _0626_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2192 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2193 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2194 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2195 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2196 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2197 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2198 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2199 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2200 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2201 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2202 VPWR net63 hold101/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2203 VGND hold101/a_285_47# hold101/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2204 net248 hold101/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2205 VGND net63 hold101/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2206 VPWR hold101/a_285_47# hold101/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2207 hold101/a_285_47# hold101/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2208 hold101/a_285_47# hold101/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2209 net248 hold101/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2210 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X2211 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X2212 VPWR acc0.A\[19\] _0609_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X2213 VGND acc0.A\[19\] _0241_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2214 _0609_/a_109_297# net46 _0241_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2215 _0241_ net46 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2216 VPWR control0.count\[1\] _0960_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2415 ps=2.83 w=0.42 l=0.15
X2217 VPWR control0.count\[2\] _0960_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2218 _0960_/a_181_47# control0.count\[0\] _0960_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0882 pd=1.26 as=0.0882 ps=1.26 w=0.42 l=0.15
X2219 VGND control0.count\[2\] _0960_/a_181_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2220 _0960_/a_27_47# control0.count\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2221 _0478_ _0960_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2222 _0478_ _0960_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2223 _0960_/a_109_47# control0.count\[1\] _0960_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2224 VPWR clknet_1_0__leaf__0457_ _0891_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X2225 _0461_ _0891_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X2226 _0461_ _0891_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X2227 VGND clknet_1_0__leaf__0457_ _0891_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X2228 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X2229 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X2230 clkload4/Y clknet_1_0__leaf__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.25
X2231 VGND clknet_1_0__leaf__0459_ clkload4/a_268_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1155 ps=1.52 w=0.55 l=0.15
X2232 clkload4/Y clknet_1_0__leaf__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.25
X2233 clkload4/Y clknet_1_0__leaf__0459_ clkload4/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0.154 pd=1.66 as=0.1155 ps=1.52 w=0.55 l=0.15
X2234 VPWR clknet_1_0__leaf__0459_ clkload4/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.25
X2235 clkload4/a_110_47# clknet_1_0__leaf__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.15
X2236 clkload4/a_268_47# clknet_1_0__leaf__0459_ clkload4/Y VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.15
X2237 VPWR clknet_1_0__leaf__0459_ clkload4/Y VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.25
X2238 VPWR acc0.A\[22\] _0222_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2239 _0222_ acc0.A\[22\] _0590_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X2240 _0590_/a_113_47# net50 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2241 _0222_ net50 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2242 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2243 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2244 VPWR clknet_1_1__leaf_clk _0857_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X2245 _0457_ _0857_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X2246 _0457_ _0857_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X2247 VGND clknet_1_1__leaf_clk _0857_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X2248 VGND _0279_ _0788_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2249 _0788_/a_68_297# _0403_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2250 _0404_ _0788_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2251 VPWR _0279_ _0788_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X2252 _0404_ _0788_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X2253 _0788_/a_150_297# _0403_ _0788_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2254 VPWR _0129_ hold16/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2255 VGND hold16/a_285_47# hold16/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2256 net163 hold16/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2257 VGND _0129_ hold16/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2258 VPWR hold16/a_285_47# hold16/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2259 hold16/a_285_47# hold16/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2260 hold16/a_285_47# hold16/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2261 net163 hold16/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2262 VPWR _0138_ hold27/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2263 VGND hold27/a_285_47# hold27/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2264 net174 hold27/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2265 VGND _0138_ hold27/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2266 VPWR hold27/a_285_47# hold27/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2267 hold27/a_285_47# hold27/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2268 hold27/a_285_47# hold27/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2269 net174 hold27/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2270 VPWR comp0.B\[3\] hold38/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2271 VGND hold38/a_285_47# hold38/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2272 net185 hold38/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2273 VGND comp0.B\[3\] hold38/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2274 VPWR hold38/a_285_47# hold38/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2275 hold38/a_285_47# hold38/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2276 hold38/a_285_47# hold38/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2277 net185 hold38/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2278 VPWR _0141_ hold49/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2279 VGND hold49/a_285_47# hold49/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2280 net196 hold49/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2281 VGND _0141_ hold49/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2282 VPWR hold49/a_285_47# hold49/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2283 hold49/a_285_47# hold49/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2284 hold49/a_285_47# hold49/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2285 net196 hold49/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2286 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2287 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2288 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2289 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2290 _0343_ control0.add VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2291 VGND control0.add _0343_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2292 _0343_ control0.add VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2293 VPWR control0.add _0343_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2294 _0642_/a_298_297# _0642_/a_27_413# _0642_/a_215_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.265 ps=2.53 w=1 l=0.15
X2295 _0642_/a_215_297# _0642_/a_27_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1359 ps=1.1 w=0.65 l=0.15
X2296 _0642_/a_298_297# _0273_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X2297 _0274_ _0642_/a_215_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.25837 ps=1.445 w=0.65 l=0.15
X2298 VPWR _0251_ _0642_/a_27_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2299 _0274_ _0642_/a_215_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2300 _0642_/a_382_47# _0252_ _0642_/a_215_297# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08775 ps=0.92 w=0.65 l=0.15
X2301 VGND _0251_ _0642_/a_27_413# VGND sky130_fd_pr__nfet_01v8 ad=0.1359 pd=1.1 as=0.1113 ps=1.37 w=0.42 l=0.15
X2302 VPWR _0252_ _0642_/a_298_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.135 ps=1.27 w=1 l=0.15
X2303 VGND _0273_ _0642_/a_382_47# VGND sky130_fd_pr__nfet_01v8 ad=0.25837 pd=1.445 as=0.091 ps=0.93 w=0.65 l=0.15
X2304 VPWR _0178_ _0573_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X2305 VGND _0573_/a_27_47# _0217_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X2306 VGND _0573_/a_27_47# _0217_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2307 _0217_ _0573_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X2308 _0217_ _0573_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2309 VGND _0178_ _0573_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X2310 VPWR _0573_/a_27_47# _0217_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2311 _0217_ _0573_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2312 _0217_ _0573_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2313 VPWR _0573_/a_27_47# _0217_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2314 net108 clknet_1_0__leaf__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2315 VGND clknet_1_0__leaf__0462_ net108 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2316 net108 clknet_1_0__leaf__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2317 VPWR clknet_1_0__leaf__0462_ net108 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2318 acc0.A\[10\] _1056_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2319 _1056_/a_891_413# _1056_/a_193_47# _1056_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2320 _1056_/a_561_413# _1056_/a_27_47# _1056_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2321 VPWR net142 _1056_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2322 acc0.A\[10\] _1056_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2323 _1056_/a_381_47# net182 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2324 VGND _1056_/a_634_159# _1056_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2325 VPWR _1056_/a_891_413# _1056_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2326 _1056_/a_466_413# _1056_/a_193_47# _1056_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2327 VPWR _1056_/a_634_159# _1056_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2328 _1056_/a_634_159# _1056_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2329 _1056_/a_634_159# _1056_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2330 _1056_/a_975_413# _1056_/a_193_47# _1056_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2331 VGND _1056_/a_1059_315# _1056_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2332 _1056_/a_193_47# _1056_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2333 _1056_/a_891_413# _1056_/a_27_47# _1056_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2334 _1056_/a_592_47# _1056_/a_193_47# _1056_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2335 VPWR _1056_/a_1059_315# _1056_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2336 _1056_/a_1017_47# _1056_/a_27_47# _1056_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2337 _1056_/a_193_47# _1056_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2338 _1056_/a_466_413# _1056_/a_27_47# _1056_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2339 VGND _1056_/a_891_413# _1056_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2340 _1056_/a_381_47# net182 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2341 VGND net142 _1056_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2342 VPWR output39/a_27_47# pp[12] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2343 pp[12] output39/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2344 VPWR net39 output39/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2345 pp[12] output39/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X2346 VGND output39/a_27_47# pp[12] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2347 VGND net39 output39/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2348 net96 clknet_1_1__leaf__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2349 VGND clknet_1_1__leaf__0460_ net96 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2350 net96 clknet_1_1__leaf__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2351 VPWR clknet_1_1__leaf__0460_ net96 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2352 VPWR net63 _0625_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2353 _0257_ _0625_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X2354 VGND net63 _0625_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2355 _0625_/a_59_75# acc0.A\[5\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2356 _0257_ _0625_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X2357 _0625_/a_145_75# acc0.A\[5\] _0625_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X2358 VGND comp0.B\[4\] _0556_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2359 _0556_/a_68_297# _0175_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2360 _0211_ _0556_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2361 VPWR comp0.B\[4\] _0556_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X2362 _0211_ _0556_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X2363 _0556_/a_150_297# _0175_ _0556_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2364 comp0.B\[7\] _1039_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2365 _1039_/a_891_413# _1039_/a_193_47# _1039_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2366 _1039_/a_561_413# _1039_/a_27_47# _1039_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2367 VPWR net125 _1039_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2368 comp0.B\[7\] _1039_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2369 _1039_/a_381_47# _0137_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2370 VGND _1039_/a_634_159# _1039_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2371 VPWR _1039_/a_891_413# _1039_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2372 _1039_/a_466_413# _1039_/a_193_47# _1039_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2373 VPWR _1039_/a_634_159# _1039_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2374 _1039_/a_634_159# _1039_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2375 _1039_/a_634_159# _1039_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2376 _1039_/a_975_413# _1039_/a_193_47# _1039_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2377 VGND _1039_/a_1059_315# _1039_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2378 _1039_/a_193_47# _1039_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2379 _1039_/a_891_413# _1039_/a_27_47# _1039_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2380 _1039_/a_592_47# _1039_/a_193_47# _1039_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2381 VPWR _1039_/a_1059_315# _1039_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2382 _1039_/a_1017_47# _1039_/a_27_47# _1039_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2383 _1039_/a_193_47# _1039_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2384 _1039_/a_466_413# _1039_/a_27_47# _1039_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2385 VGND _1039_/a_891_413# _1039_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2386 _1039_/a_381_47# _0137_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2387 VGND net125 _1039_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2388 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X2389 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X2390 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2391 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2392 _0240_ net44 _0608_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.348 pd=2.78 as=0.21 ps=2.42 w=1 l=0.15
X2393 VPWR _0239_ _0240_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.7 l=0.15
X2394 _0608_/a_27_47# net44 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X2395 _0240_ _0239_ _0608_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2396 _0608_/a_109_297# acc0.A\[17\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2397 VGND acc0.A\[17\] _0608_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2398 VGND comp0.B\[12\] _0539_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2399 _0539_/a_68_297# _0176_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2400 _0202_ _0539_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2401 VPWR comp0.B\[12\] _0539_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X2402 _0202_ _0539_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X2403 _0539_/a_150_297# _0176_ _0539_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2404 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2405 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2406 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2407 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2408 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2409 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2410 net147 clknet_1_0__leaf__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2411 VGND clknet_1_0__leaf__0465_ net147 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2412 net147 clknet_1_0__leaf__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2413 VPWR clknet_1_0__leaf__0465_ net147 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2414 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2415 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2416 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X2417 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X2418 control0.count\[3\] _1072_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2419 _1072_/a_891_413# _1072_/a_193_47# _1072_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2420 _1072_/a_561_413# _1072_/a_27_47# _1072_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2421 VPWR clknet_1_0__leaf_clk _1072_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2422 control0.count\[3\] _1072_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2423 _1072_/a_381_47# _0170_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2424 VGND _1072_/a_634_159# _1072_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2425 VPWR _1072_/a_891_413# _1072_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2426 _1072_/a_466_413# _1072_/a_193_47# _1072_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2427 VPWR _1072_/a_634_159# _1072_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2428 _1072_/a_634_159# _1072_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2429 _1072_/a_634_159# _1072_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2430 _1072_/a_975_413# _1072_/a_193_47# _1072_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2431 VGND _1072_/a_1059_315# _1072_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2432 _1072_/a_193_47# _1072_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2433 _1072_/a_891_413# _1072_/a_27_47# _1072_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2434 _1072_/a_592_47# _1072_/a_193_47# _1072_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2435 VPWR _1072_/a_1059_315# _1072_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2436 _1072_/a_1017_47# _1072_/a_27_47# _1072_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2437 _1072_/a_193_47# _1072_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2438 _1072_/a_466_413# _1072_/a_27_47# _1072_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2439 VGND _1072_/a_891_413# _1072_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2440 _1072_/a_381_47# _0170_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2441 VGND clknet_1_0__leaf_clk _1072_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2442 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2443 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2444 VPWR _0787_/a_80_21# _0403_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X2445 _0787_/a_209_297# _0402_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.65 pd=5.3 as=0 ps=0 w=1 l=0.15
X2446 _0787_/a_303_47# _0285_ _0787_/a_209_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.208 ps=1.94 w=0.65 l=0.15
X2447 _0787_/a_209_47# _0402_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2448 VGND _0787_/a_80_21# _0403_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.17225 ps=1.83 w=0.65 l=0.15
X2449 VGND _0284_ _0787_/a_80_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2145 ps=1.96 w=0.65 l=0.15
X2450 _0787_/a_80_21# _0281_ _0787_/a_303_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2451 VPWR _0285_ _0787_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2452 _0787_/a_80_21# _0284_ _0787_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0 ps=0 w=1 l=0.15
X2453 _0787_/a_209_297# _0281_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2454 VGND _0346_ _0856_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X2455 _0856_/a_510_47# _0456_ _0856_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X2456 _0856_/a_79_21# _0345_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X2457 VPWR _0456_ _0856_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2458 _0856_/a_79_21# _0264_ _0856_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X2459 _0856_/a_297_297# _0346_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2460 _0856_/a_79_21# _0345_ _0856_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X2461 VPWR _0856_/a_79_21# _0080_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2462 VGND _0856_/a_79_21# _0080_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2463 _0856_/a_215_47# _0264_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2464 VPWR control0.count\[2\] hold17/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2465 VGND hold17/a_285_47# hold17/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2466 net164 hold17/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2467 VGND control0.count\[2\] hold17/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2468 VPWR hold17/a_285_47# hold17/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2469 hold17/a_285_47# hold17/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2470 hold17/a_285_47# hold17/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2471 net164 hold17/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2472 VPWR acc0.A\[2\] hold28/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2473 VGND hold28/a_285_47# hold28/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2474 net175 hold28/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2475 VGND acc0.A\[2\] hold28/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2476 VPWR hold28/a_285_47# hold28/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2477 hold28/a_285_47# hold28/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2478 hold28/a_285_47# hold28/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2479 net175 hold28/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2480 VPWR _0132_ hold39/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2481 VGND hold39/a_285_47# hold39/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2482 net186 hold39/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2483 VGND _0132_ hold39/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2484 VPWR hold39/a_285_47# hold39/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2485 hold39/a_285_47# hold39/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2486 hold39/a_285_47# hold39/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2487 net186 hold39/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2488 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X2489 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X2490 _0342_ _0340_ _0710_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
X2491 _0342_ _0340_ _0710_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2492 VPWR _0339_ _0710_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.135 ps=1.27 w=1 l=0.15
X2493 _0710_/a_109_297# _0220_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2494 _0710_/a_381_47# _0220_ _0342_ VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.169 ps=1.82 w=0.65 l=0.15
X2495 _0710_/a_109_297# _0341_ _0342_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2496 _0710_/a_109_47# _0341_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X2497 VGND _0339_ _0710_/a_381_47# VGND sky130_fd_pr__nfet_01v8 ad=0.234 pd=2.02 as=0.06825 ps=0.86 w=0.65 l=0.15
X2498 VPWR acc0.A\[6\] _0273_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2499 _0273_ acc0.A\[6\] _0641_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X2500 _0641_/a_113_47# net64 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2501 _0273_ net64 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2502 VPWR _0216_ _0572_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X2503 _0572_/a_27_297# _0195_ _0572_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X2504 VGND _0216_ _0572_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X2505 _0124_ _0572_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2506 _0572_/a_27_297# _0195_ _0572_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X2507 _0572_/a_109_297# net155 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2508 _0572_/a_373_47# net155 _0572_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2509 _0124_ _0572_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2510 _0572_/a_109_297# net210 _0572_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2511 _0572_/a_109_47# net210 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2512 acc0.A\[9\] _1055_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2513 _1055_/a_891_413# _1055_/a_193_47# _1055_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2514 _1055_/a_561_413# _1055_/a_27_47# _1055_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2515 VPWR net141 _1055_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2516 acc0.A\[9\] _1055_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2517 _1055_/a_381_47# net179 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2518 VGND _1055_/a_634_159# _1055_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2519 VPWR _1055_/a_891_413# _1055_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2520 _1055_/a_466_413# _1055_/a_193_47# _1055_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2521 VPWR _1055_/a_634_159# _1055_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2522 _1055_/a_634_159# _1055_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2523 _1055_/a_634_159# _1055_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2524 _1055_/a_975_413# _1055_/a_193_47# _1055_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2525 VGND _1055_/a_1059_315# _1055_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2526 _1055_/a_193_47# _1055_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2527 _1055_/a_891_413# _1055_/a_27_47# _1055_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2528 _1055_/a_592_47# _1055_/a_193_47# _1055_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2529 VPWR _1055_/a_1059_315# _1055_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2530 _1055_/a_1017_47# _1055_/a_27_47# _1055_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2531 _1055_/a_193_47# _1055_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2532 _1055_/a_466_413# _1055_/a_27_47# _1055_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2533 VGND _1055_/a_891_413# _1055_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2534 _1055_/a_381_47# net179 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2535 VGND net141 _1055_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2536 VPWR _0432_ _0839_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X2537 VGND _0432_ _0444_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2538 _0839_/a_109_297# _0443_ _0444_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2539 _0444_ _0443_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2540 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2541 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2542 VPWR net62 _0624_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2543 _0256_ _0624_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X2544 VGND net62 _0624_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2545 _0624_/a_59_75# acc0.A\[4\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2546 _0256_ _0624_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X2547 _0624_/a_145_75# acc0.A\[4\] _0624_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X2548 _0555_/a_240_47# net28 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X2549 _0135_ _0555_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X2550 VGND _0208_ _0555_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2551 _0555_/a_51_297# net204 _0555_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X2552 _0555_/a_149_47# _0210_ _0555_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X2553 _0555_/a_240_47# _0173_ _0555_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2554 VPWR _0208_ _0555_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X2555 _0135_ _0555_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X2556 _0555_/a_149_47# net204 _0555_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2557 _0555_/a_245_297# _0173_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2558 VPWR _0210_ _0555_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2559 _0555_/a_512_297# net28 _0555_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2560 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2561 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2562 comp0.B\[6\] _1038_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2563 _1038_/a_891_413# _1038_/a_193_47# _1038_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2564 _1038_/a_561_413# _1038_/a_27_47# _1038_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2565 VPWR net124 _1038_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2566 comp0.B\[6\] _1038_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2567 _1038_/a_381_47# net172 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2568 VGND _1038_/a_634_159# _1038_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2569 VPWR _1038_/a_891_413# _1038_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2570 _1038_/a_466_413# _1038_/a_193_47# _1038_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2571 VPWR _1038_/a_634_159# _1038_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2572 _1038_/a_634_159# _1038_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2573 _1038_/a_634_159# _1038_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2574 _1038_/a_975_413# _1038_/a_193_47# _1038_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2575 VGND _1038_/a_1059_315# _1038_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2576 _1038_/a_193_47# _1038_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2577 _1038_/a_891_413# _1038_/a_27_47# _1038_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2578 _1038_/a_592_47# _1038_/a_193_47# _1038_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2579 VPWR _1038_/a_1059_315# _1038_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2580 _1038_/a_1017_47# _1038_/a_27_47# _1038_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2581 _1038_/a_193_47# _1038_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2582 _1038_/a_466_413# _1038_/a_27_47# _1038_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2583 VGND _1038_/a_891_413# _1038_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2584 _1038_/a_381_47# net172 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2585 VGND net124 _1038_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2586 net100 clknet_1_0__leaf__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2587 VGND clknet_1_0__leaf__0461_ net100 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2588 net100 clknet_1_0__leaf__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2589 VPWR clknet_1_0__leaf__0461_ net100 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2590 _0538_/a_240_47# net21 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X2591 _0143_ _0538_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X2592 VGND _0172_ _0538_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2593 _0538_/a_51_297# net183 _0538_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X2594 _0538_/a_149_47# _0201_ _0538_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X2595 _0538_/a_240_47# _0174_ _0538_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2596 VPWR _0172_ _0538_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X2597 _0143_ _0538_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X2598 _0538_/a_149_47# net183 _0538_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2599 _0538_/a_245_297# _0174_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2600 VPWR _0201_ _0538_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2601 _0538_/a_512_297# net21 _0538_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2602 VPWR net44 _0607_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X2603 _0607_/a_27_297# net43 _0607_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X2604 VGND net44 _0607_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X2605 _0239_ _0607_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2606 _0607_/a_27_297# net43 _0607_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X2607 _0607_/a_109_297# acc0.A\[17\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2608 _0607_/a_373_47# acc0.A\[17\] _0607_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2609 _0239_ _0607_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2610 _0607_/a_109_297# acc0.A\[16\] _0607_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2611 _0607_/a_109_47# acc0.A\[16\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2612 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2613 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2614 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2615 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2616 net81 clknet_1_1__leaf__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2617 VGND clknet_1_1__leaf__0459_ net81 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2618 net81 clknet_1_1__leaf__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2619 VPWR clknet_1_1__leaf__0459_ net81 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2620 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X2621 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X2622 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X2623 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X2624 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2625 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2626 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2627 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2628 control0.count\[2\] _1071_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2629 _1071_/a_891_413# _1071_/a_193_47# _1071_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2630 _1071_/a_561_413# _1071_/a_27_47# _1071_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2631 VPWR clknet_1_0__leaf_clk _1071_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2632 control0.count\[2\] _1071_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2633 _1071_/a_381_47# _0169_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2634 VGND _1071_/a_634_159# _1071_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2635 VPWR _1071_/a_891_413# _1071_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2636 _1071_/a_466_413# _1071_/a_193_47# _1071_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2637 VPWR _1071_/a_634_159# _1071_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2638 _1071_/a_634_159# _1071_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2639 _1071_/a_634_159# _1071_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2640 _1071_/a_975_413# _1071_/a_193_47# _1071_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2641 VGND _1071_/a_1059_315# _1071_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2642 _1071_/a_193_47# _1071_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2643 _1071_/a_891_413# _1071_/a_27_47# _1071_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2644 _1071_/a_592_47# _1071_/a_193_47# _1071_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2645 VPWR _1071_/a_1059_315# _1071_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2646 _1071_/a_1017_47# _1071_/a_27_47# _1071_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2647 _1071_/a_193_47# _1071_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2648 _1071_/a_466_413# _1071_/a_27_47# _1071_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2649 VGND _1071_/a_891_413# _1071_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2650 _1071_/a_381_47# _0169_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2651 VGND clknet_1_0__leaf_clk _1071_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2652 VPWR clknet_1_1__leaf__0457_ _0924_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X2653 _0464_ _0924_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X2654 _0464_ _0924_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X2655 VGND clknet_1_1__leaf__0457_ _0924_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X2656 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2657 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2658 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2659 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2660 _0855_/a_81_21# net234 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X2661 _0855_/a_299_297# net234 _0855_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X2662 VPWR _0855_/a_81_21# _0456_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2663 VPWR net149 _0855_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2664 VGND _0855_/a_81_21# _0456_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2665 VGND _0350_ _0855_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X2666 _0855_/a_299_297# _0350_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2667 _0855_/a_384_47# net149 _0855_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2668 VPWR _0786_/a_80_21# _0402_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X2669 _0786_/a_80_21# _0289_ _0786_/a_472_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.31 ps=2.62 w=1 l=0.15
X2670 VPWR _0401_ _0786_/a_217_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.545 ps=5.09 w=1 l=0.15
X2671 VGND _0283_ _0786_/a_80_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.35425 ps=3.69 w=0.65 l=0.15
X2672 VGND _0786_/a_80_21# _0402_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.17225 ps=1.83 w=0.65 l=0.15
X2673 _0786_/a_300_47# _0401_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X2674 _0786_/a_217_297# _0295_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2675 _0786_/a_80_21# _0295_ _0786_/a_300_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2676 _0786_/a_472_297# _0283_ _0786_/a_217_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2677 _0786_/a_80_21# _0289_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2678 VPWR acc0.A\[15\] hold18/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2679 VGND hold18/a_285_47# hold18/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2680 net165 hold18/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2681 VGND acc0.A\[15\] hold18/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2682 VPWR hold18/a_285_47# hold18/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2683 hold18/a_285_47# hold18/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2684 hold18/a_285_47# hold18/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2685 net165 hold18/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2686 VPWR acc0.A\[22\] hold29/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2687 VGND hold29/a_285_47# hold29/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2688 net176 hold29/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2689 VGND acc0.A\[22\] hold29/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2690 VPWR hold29/a_285_47# hold29/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2691 hold29/a_285_47# hold29/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2692 hold29/a_285_47# hold29/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2693 net176 hold29/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2694 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2695 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2696 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X2697 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X2698 _0272_ _0640_/a_215_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X2699 _0640_/a_109_53# _0271_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2700 _0640_/a_215_297# _0640_/a_109_53# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X2701 _0272_ _0640_/a_215_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.10187 ps=0.99 w=0.65 l=0.15
X2702 _0640_/a_392_297# _0255_ _0640_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.04515 pd=0.635 as=0.06825 ps=0.745 w=0.42 l=0.15
X2703 _0640_/a_465_297# _0257_ _0640_/a_392_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.04515 ps=0.635 w=0.42 l=0.15
X2704 _0640_/a_215_297# _0257_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2705 VPWR _0254_ _0640_/a_465_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06405 ps=0.725 w=0.42 l=0.15
X2706 _0640_/a_297_297# _0640_/a_109_53# _0640_/a_215_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X2707 _0640_/a_109_53# _0271_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2708 VGND _0255_ _0640_/a_215_297# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X2709 VGND _0254_ _0640_/a_215_297# VGND sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X2710 VPWR _0216_ _0571_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X2711 _0571_/a_27_297# _0195_ _0571_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X2712 VGND _0216_ _0571_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X2713 _0125_ _0571_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2714 _0571_/a_27_297# _0195_ _0571_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X2715 _0571_/a_109_297# acc0.A\[27\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2716 _0571_/a_373_47# acc0.A\[27\] _0571_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2717 _0125_ _0571_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2718 _0571_/a_109_297# net155 _0571_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2719 _0571_/a_109_47# net155 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2720 acc0.A\[8\] _1054_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2721 _1054_/a_891_413# _1054_/a_193_47# _1054_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2722 _1054_/a_561_413# _1054_/a_27_47# _1054_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2723 VPWR net140 _1054_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2724 acc0.A\[8\] _1054_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2725 _1054_/a_381_47# net169 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2726 VGND _1054_/a_634_159# _1054_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2727 VPWR _1054_/a_891_413# _1054_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2728 _1054_/a_466_413# _1054_/a_193_47# _1054_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2729 VPWR _1054_/a_634_159# _1054_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2730 _1054_/a_634_159# _1054_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2731 _1054_/a_634_159# _1054_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2732 _1054_/a_975_413# _1054_/a_193_47# _1054_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2733 VGND _1054_/a_1059_315# _1054_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2734 _1054_/a_193_47# _1054_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2735 _1054_/a_891_413# _1054_/a_27_47# _1054_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2736 _1054_/a_592_47# _1054_/a_193_47# _1054_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2737 VPWR _1054_/a_1059_315# _1054_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2738 _1054_/a_1017_47# _1054_/a_27_47# _1054_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2739 _1054_/a_193_47# _1054_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2740 _1054_/a_466_413# _1054_/a_27_47# _1054_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2741 VGND _1054_/a_891_413# _1054_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2742 _1054_/a_381_47# net169 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2743 VGND net140 _1054_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2744 _0769_/a_81_21# _0244_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X2745 _0769_/a_299_297# _0244_ _0769_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X2746 VPWR _0769_/a_81_21# _0389_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2747 VPWR _0386_ _0769_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2748 VGND _0769_/a_81_21# _0389_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2749 VGND _0388_ _0769_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X2750 _0769_/a_299_297# _0388_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2751 _0769_/a_384_47# _0386_ _0769_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2752 VPWR _0431_ _0838_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X2753 VGND _0431_ _0443_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2754 _0838_/a_109_297# _0271_ _0443_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2755 _0443_ _0271_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2756 VPWR acc0.A\[5\] _0623_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X2757 VGND acc0.A\[5\] _0255_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2758 _0623_/a_109_297# net63 _0255_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2759 _0255_ net63 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2760 VGND net160 _0554_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2761 _0554_/a_68_297# _0175_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2762 _0210_ _0554_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2763 VPWR net160 _0554_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X2764 _0210_ _0554_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X2765 _0554_/a_150_297# _0175_ _0554_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2766 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X2767 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X2768 comp0.B\[5\] _1037_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2769 _1037_/a_891_413# _1037_/a_193_47# _1037_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2770 _1037_/a_561_413# _1037_/a_27_47# _1037_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2771 VPWR net123 _1037_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2772 comp0.B\[5\] _1037_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2773 _1037_/a_381_47# _0135_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2774 VGND _1037_/a_634_159# _1037_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2775 VPWR _1037_/a_891_413# _1037_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2776 _1037_/a_466_413# _1037_/a_193_47# _1037_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2777 VPWR _1037_/a_634_159# _1037_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2778 _1037_/a_634_159# _1037_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2779 _1037_/a_634_159# _1037_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2780 _1037_/a_975_413# _1037_/a_193_47# _1037_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2781 VGND _1037_/a_1059_315# _1037_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2782 _1037_/a_193_47# _1037_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2783 _1037_/a_891_413# _1037_/a_27_47# _1037_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2784 _1037_/a_592_47# _1037_/a_193_47# _1037_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2785 VPWR _1037_/a_1059_315# _1037_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2786 _1037_/a_1017_47# _1037_/a_27_47# _1037_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2787 _1037_/a_193_47# _1037_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2788 _1037_/a_466_413# _1037_/a_27_47# _1037_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2789 VGND _1037_/a_891_413# _1037_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2790 _1037_/a_381_47# _0135_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2791 VGND net123 _1037_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2792 net87 clknet_1_0__leaf__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2793 VGND clknet_1_0__leaf__0459_ net87 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2794 net87 clknet_1_0__leaf__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2795 VPWR clknet_1_0__leaf__0459_ net87 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2796 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2797 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2798 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2799 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2800 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2801 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2802 _0238_ _0606_/a_215_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0 ps=0 w=1 l=0.15
X2803 _0606_/a_109_53# _0237_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2804 _0606_/a_215_297# _0606_/a_109_53# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2415 pd=2.83 as=0 ps=0 w=0.42 l=0.15
X2805 _0238_ _0606_/a_215_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X2806 _0606_/a_392_297# _0236_ _0606_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0903 pd=1.27 as=0.1365 ps=1.49 w=0.42 l=0.15
X2807 _0606_/a_465_297# _0234_ _0606_/a_392_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1281 pd=1.45 as=0 ps=0 w=0.42 l=0.15
X2808 _0606_/a_215_297# _0234_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2809 VPWR _0225_ _0606_/a_465_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2810 _0606_/a_297_297# _0606_/a_109_53# _0606_/a_215_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2811 _0606_/a_109_53# _0237_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2812 VGND _0236_ _0606_/a_215_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2813 VGND _0225_ _0606_/a_215_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2814 VGND comp0.B\[13\] _0537_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2815 _0537_/a_68_297# _0176_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2816 _0201_ _0537_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2817 VPWR comp0.B\[13\] _0537_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X2818 _0201_ _0537_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X2819 _0537_/a_150_297# _0176_ _0537_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2820 net76 clknet_1_1__leaf__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2821 VGND clknet_1_1__leaf__0458_ net76 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2822 net76 clknet_1_1__leaf__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2823 VPWR clknet_1_1__leaf__0458_ net76 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2824 net138 clknet_1_0__leaf__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2825 VGND clknet_1_0__leaf__0465_ net138 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2826 net138 clknet_1_0__leaf__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2827 VPWR clknet_1_0__leaf__0465_ net138 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2828 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2829 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2830 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X2831 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X2832 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2833 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2834 net119 clknet_1_1__leaf__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2835 VGND clknet_1_1__leaf__0463_ net119 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2836 net119 clknet_1_1__leaf__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2837 VPWR clknet_1_1__leaf__0463_ net119 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2838 control0.count\[1\] _1070_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2839 _1070_/a_891_413# _1070_/a_193_47# _1070_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2840 _1070_/a_561_413# _1070_/a_27_47# _1070_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2841 VPWR clknet_1_0__leaf_clk _1070_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2842 control0.count\[1\] _1070_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2843 _1070_/a_381_47# _0168_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2844 VGND _1070_/a_634_159# _1070_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2845 VPWR _1070_/a_891_413# _1070_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2846 _1070_/a_466_413# _1070_/a_193_47# _1070_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2847 VPWR _1070_/a_634_159# _1070_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2848 _1070_/a_634_159# _1070_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2849 _1070_/a_634_159# _1070_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2850 _1070_/a_975_413# _1070_/a_193_47# _1070_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2851 VGND _1070_/a_1059_315# _1070_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2852 _1070_/a_193_47# _1070_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2853 _1070_/a_891_413# _1070_/a_27_47# _1070_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2854 _1070_/a_592_47# _1070_/a_193_47# _1070_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2855 VPWR _1070_/a_1059_315# _1070_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2856 _1070_/a_1017_47# _1070_/a_27_47# _1070_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2857 _1070_/a_193_47# _1070_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2858 _1070_/a_466_413# _1070_/a_27_47# _1070_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2859 VGND _1070_/a_891_413# _1070_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2860 _1070_/a_381_47# _0168_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2861 VGND clknet_1_0__leaf_clk _1070_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2862 net133 clknet_1_0__leaf__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X2863 VGND clknet_1_0__leaf__0464_ net133 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X2864 net133 clknet_1_0__leaf__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2865 VPWR clknet_1_0__leaf__0464_ net133 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2866 VGND _0347_ _0854_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X2867 _0854_/a_510_47# _0455_ _0854_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X2868 _0854_/a_79_21# _0399_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X2869 VPWR _0455_ _0854_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2870 _0854_/a_79_21# _0454_ _0854_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X2871 _0854_/a_297_297# _0347_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2872 _0854_/a_79_21# _0399_ _0854_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X2873 VPWR _0854_/a_79_21# _0081_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2874 VGND _0854_/a_79_21# _0081_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2875 _0854_/a_215_47# _0454_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2876 _0785_/a_81_21# _0292_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X2877 _0785_/a_299_297# _0292_ _0785_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X2878 VPWR _0785_/a_81_21# _0401_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X2879 VPWR _0259_ _0785_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2880 VGND _0785_/a_81_21# _0401_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2881 VGND _0275_ _0785_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X2882 _0785_/a_299_297# _0275_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2883 _0785_/a_384_47# _0259_ _0785_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2884 VPWR _0114_ hold19/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2885 VGND hold19/a_285_47# hold19/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2886 net166 hold19/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2887 VGND _0114_ hold19/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2888 VPWR hold19/a_285_47# hold19/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X2889 hold19/a_285_47# hold19/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2890 hold19/a_285_47# hold19/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X2891 net166 hold19/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2892 VPWR _0216_ _0570_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X2893 _0570_/a_27_297# _0195_ _0570_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X2894 VGND _0216_ _0570_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X2895 _0126_ _0570_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2896 _0570_/a_27_297# _0195_ _0570_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X2897 _0570_/a_109_297# net190 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2898 _0570_/a_373_47# net190 _0570_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2899 _0126_ _0570_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2900 _0570_/a_109_297# net197 _0570_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2901 _0570_/a_109_47# net197 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2902 acc0.A\[7\] _1053_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2903 _1053_/a_891_413# _1053_/a_193_47# _1053_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2904 _1053_/a_561_413# _1053_/a_27_47# _1053_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2905 VPWR net139 _1053_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2906 acc0.A\[7\] _1053_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2907 _1053_/a_381_47# _0151_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2908 VGND _1053_/a_634_159# _1053_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2909 VPWR _1053_/a_891_413# _1053_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2910 _1053_/a_466_413# _1053_/a_193_47# _1053_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2911 VPWR _1053_/a_634_159# _1053_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2912 _1053_/a_634_159# _1053_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2913 _1053_/a_634_159# _1053_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2914 _1053_/a_975_413# _1053_/a_193_47# _1053_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2915 VGND _1053_/a_1059_315# _1053_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2916 _1053_/a_193_47# _1053_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2917 _1053_/a_891_413# _1053_/a_27_47# _1053_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2918 _1053_/a_592_47# _1053_/a_193_47# _1053_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2919 VPWR _1053_/a_1059_315# _1053_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2920 _1053_/a_1017_47# _1053_/a_27_47# _1053_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2921 _1053_/a_193_47# _1053_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2922 _1053_/a_466_413# _1053_/a_27_47# _1053_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2923 VGND _1053_/a_891_413# _1053_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2924 _1053_/a_381_47# _0151_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2925 VGND net139 _1053_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2926 _0837_/a_585_47# _0442_ _0837_/a_266_47# VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.11863 ps=1.015 w=0.65 l=0.15
X2927 VGND _0440_ _0837_/a_266_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.07 as=0.117 ps=1.01 w=0.65 l=0.15
X2928 VPWR _0837_/a_81_21# _0085_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3125 pd=1.625 as=0.26 ps=2.52 w=1 l=0.15
X2929 _0837_/a_81_21# _0172_ _0837_/a_585_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X2930 VGND _0837_/a_81_21# _0085_ VGND sky130_fd_pr__nfet_01v8 ad=0.20312 pd=1.275 as=0.169 ps=1.82 w=0.65 l=0.15
X2931 _0837_/a_266_297# _0346_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.3125 ps=1.625 w=1 l=0.15
X2932 _0837_/a_368_297# _0440_ _0837_/a_266_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=1.42 as=0.18 ps=1.36 w=1 l=0.15
X2933 _0837_/a_266_47# _0441_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.11863 pd=1.015 as=0.1365 ps=1.07 w=0.65 l=0.15
X2934 _0837_/a_266_47# _0346_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.20312 ps=1.275 w=0.65 l=0.15
X2935 _0837_/a_81_21# _0441_ _0837_/a_368_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.21 ps=1.42 w=1 l=0.15
X2936 _0837_/a_81_21# _0172_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.15 ps=1.3 w=1 l=0.15
X2937 VPWR _0442_ _0837_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.15 pd=1.3 as=0.1375 ps=1.275 w=1 l=0.15
X2938 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X2939 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X2940 _0388_ _0310_ _0768_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.348 pd=2.78 as=0.21 ps=2.42 w=1 l=0.15
X2941 VPWR _0240_ _0388_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.7 l=0.15
X2942 _0768_/a_27_47# _0310_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X2943 _0388_ _0240_ _0768_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2944 _0768_/a_109_297# _0387_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2945 VGND _0387_ _0768_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2946 VGND acc0.A\[28\] _0699_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X2947 _0699_/a_68_297# net56 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2948 _0331_ _0699_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2949 VPWR acc0.A\[28\] _0699_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X2950 _0331_ _0699_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X2951 _0699_/a_150_297# net56 _0699_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2952 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X2953 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X2954 VPWR _0252_ _0254_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X2955 _0254_ _0251_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.165 ps=1.33 w=1 l=0.15
X2956 _0622_/a_193_47# _0252_ _0622_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X2957 _0254_ _0251_ _0622_/a_193_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10725 ps=0.98 w=0.65 l=0.15
X2958 _0254_ _0253_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2959 _0622_/a_109_47# _0253_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2960 _0553_/a_240_47# net29 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X2961 _0136_ _0553_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X2962 VGND _0208_ _0553_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2963 _0553_/a_51_297# net171 _0553_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X2964 _0553_/a_149_47# _0209_ _0553_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X2965 _0553_/a_240_47# _0174_ _0553_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2966 VPWR _0208_ _0553_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X2967 _0136_ _0553_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X2968 _0553_/a_149_47# net171 _0553_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X2969 _0553_/a_245_297# _0174_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2970 VPWR _0209_ _0553_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2971 _0553_/a_512_297# net29 _0553_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X2972 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X2973 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X2974 comp0.B\[4\] _1036_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X2975 _1036_/a_891_413# _1036_/a_193_47# _1036_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X2976 _1036_/a_561_413# _1036_/a_27_47# _1036_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X2977 VPWR net122 _1036_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X2978 comp0.B\[4\] _1036_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X2979 _1036_/a_381_47# net161 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X2980 VGND _1036_/a_634_159# _1036_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X2981 VPWR _1036_/a_891_413# _1036_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X2982 _1036_/a_466_413# _1036_/a_193_47# _1036_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2983 VPWR _1036_/a_634_159# _1036_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2984 _1036_/a_634_159# _1036_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X2985 _1036_/a_634_159# _1036_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X2986 _1036_/a_975_413# _1036_/a_193_47# _1036_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X2987 VGND _1036_/a_1059_315# _1036_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X2988 _1036_/a_193_47# _1036_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X2989 _1036_/a_891_413# _1036_/a_27_47# _1036_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2990 _1036_/a_592_47# _1036_/a_193_47# _1036_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X2991 VPWR _1036_/a_1059_315# _1036_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2992 _1036_/a_1017_47# _1036_/a_27_47# _1036_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X2993 _1036_/a_193_47# _1036_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X2994 _1036_/a_466_413# _1036_/a_27_47# _1036_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X2995 VGND _1036_/a_891_413# _1036_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X2996 _1036_/a_381_47# net161 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X2997 VGND net122 _1036_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X2998 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X2999 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X3000 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3001 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3002 _0536_/a_240_47# net22 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X3003 _0144_ _0536_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X3004 VGND _0172_ _0536_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3005 _0536_/a_51_297# net157 _0536_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X3006 _0536_/a_149_47# _0200_ _0536_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X3007 _0536_/a_240_47# _0174_ _0536_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3008 VPWR _0172_ _0536_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X3009 _0144_ _0536_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X3010 _0536_/a_149_47# net157 _0536_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3011 _0536_/a_245_297# _0174_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3012 VPWR _0200_ _0536_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3013 _0536_/a_512_297# net22 _0536_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3014 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3015 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3016 VPWR _0228_ _0605_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X3017 VGND _0228_ _0237_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X3018 _0605_/a_109_297# _0227_ _0237_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X3019 _0237_ _0227_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3020 acc0.A\[19\] _1019_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3021 _1019_/a_891_413# _1019_/a_193_47# _1019_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3022 _1019_/a_561_413# _1019_/a_27_47# _1019_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3023 VPWR net105 _1019_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3024 acc0.A\[19\] _1019_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3025 _1019_/a_381_47# net207 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3026 VGND _1019_/a_634_159# _1019_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3027 VPWR _1019_/a_891_413# _1019_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3028 _1019_/a_466_413# _1019_/a_193_47# _1019_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3029 VPWR _1019_/a_634_159# _1019_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3030 _1019_/a_634_159# _1019_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3031 _1019_/a_634_159# _1019_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3032 _1019_/a_975_413# _1019_/a_193_47# _1019_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3033 VGND _1019_/a_1059_315# _1019_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3034 _1019_/a_193_47# _1019_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3035 _1019_/a_891_413# _1019_/a_27_47# _1019_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3036 _1019_/a_592_47# _1019_/a_193_47# _1019_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3037 VPWR _1019_/a_1059_315# _1019_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3038 _1019_/a_1017_47# _1019_/a_27_47# _1019_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3039 _1019_/a_193_47# _1019_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3040 _1019_/a_466_413# _1019_/a_27_47# _1019_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3041 VGND _1019_/a_891_413# _1019_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3042 _1019_/a_381_47# net207 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3043 VGND net105 _1019_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3044 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X3045 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X3046 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X3047 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X3048 VPWR clknet_0__0465_ clkbuf_1_1__f__0465_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X3049 VPWR clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X3050 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3051 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3052 VPWR clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3053 VPWR clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3054 clkbuf_1_1__f__0465_/a_110_47# clknet_0__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3055 clkbuf_1_1__f__0465_/a_110_47# clknet_0__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X3056 VGND clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X3057 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3058 VGND clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3059 clkbuf_1_1__f__0465_/a_110_47# clknet_0__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3060 VGND clknet_0__0465_ clkbuf_1_1__f__0465_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3061 VGND clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3062 VPWR clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3063 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3064 VGND clknet_0__0465_ clkbuf_1_1__f__0465_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3065 VGND clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3066 VPWR clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3067 VGND clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3068 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3069 clkbuf_1_1__f__0465_/a_110_47# clknet_0__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3070 VPWR clknet_0__0465_ clkbuf_1_1__f__0465_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3071 VPWR clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3072 VPWR clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3073 VGND clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3074 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3075 VGND clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3076 VGND clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3077 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3078 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3079 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3080 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3081 VPWR clkbuf_1_1__f__0465_/a_110_47# clknet_1_1__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3082 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3083 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3084 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3085 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3086 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3087 clknet_1_1__leaf__0465_ clkbuf_1_1__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3088 _0519_/a_81_21# _0191_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X3089 _0519_/a_299_297# _0191_ _0519_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X3090 VPWR _0519_/a_81_21# _0152_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X3091 VPWR net168 _0519_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3092 VGND _0519_/a_81_21# _0152_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3093 VGND _0179_ _0519_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X3094 _0519_/a_299_297# _0179_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3095 _0519_/a_384_47# net168 _0519_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3096 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3097 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3098 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X3099 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X3100 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3101 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3102 net44 _0999_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3103 _0999_/a_891_413# _0999_/a_193_47# _0999_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3104 _0999_/a_561_413# _0999_/a_27_47# _0999_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3105 VPWR net85 _0999_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3106 net44 _0999_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3107 _0999_/a_381_47# _0097_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3108 VGND _0999_/a_634_159# _0999_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3109 VPWR _0999_/a_891_413# _0999_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3110 _0999_/a_466_413# _0999_/a_193_47# _0999_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3111 VPWR _0999_/a_634_159# _0999_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3112 _0999_/a_634_159# _0999_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3113 _0999_/a_634_159# _0999_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3114 _0999_/a_975_413# _0999_/a_193_47# _0999_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3115 VGND _0999_/a_1059_315# _0999_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3116 _0999_/a_193_47# _0999_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3117 _0999_/a_891_413# _0999_/a_27_47# _0999_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3118 _0999_/a_592_47# _0999_/a_193_47# _0999_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3119 VPWR _0999_/a_1059_315# _0999_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3120 _0999_/a_1017_47# _0999_/a_27_47# _0999_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3121 _0999_/a_193_47# _0999_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3122 _0999_/a_466_413# _0999_/a_27_47# _0999_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3123 VGND _0999_/a_891_413# _0999_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3124 _0999_/a_381_47# _0097_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3125 VGND net85 _0999_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3126 VGND _0218_ _0853_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X3127 _0853_/a_68_297# net47 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3128 _0455_ _0853_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3129 VPWR _0218_ _0853_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X3130 _0455_ _0853_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X3131 _0853_/a_150_297# net47 _0853_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3132 VPWR acc0.A\[14\] _0400_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3133 _0400_ acc0.A\[14\] _0784_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X3134 _0784_/a_113_47# net41 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3135 _0400_ net41 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3136 VPWR A[0] input1/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X3137 net1 input1/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X3138 net1 input1/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X3139 VGND A[0] input1/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X3140 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X3141 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X3142 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3143 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3144 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X3145 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X3146 acc0.A\[6\] _1052_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3147 _1052_/a_891_413# _1052_/a_193_47# _1052_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3148 _1052_/a_561_413# _1052_/a_27_47# _1052_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3149 VPWR net138 _1052_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3150 acc0.A\[6\] _1052_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3151 _1052_/a_381_47# _0150_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3152 VGND _1052_/a_634_159# _1052_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3153 VPWR _1052_/a_891_413# _1052_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3154 _1052_/a_466_413# _1052_/a_193_47# _1052_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3155 VPWR _1052_/a_634_159# _1052_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3156 _1052_/a_634_159# _1052_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3157 _1052_/a_634_159# _1052_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3158 _1052_/a_975_413# _1052_/a_193_47# _1052_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3159 VGND _1052_/a_1059_315# _1052_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3160 _1052_/a_193_47# _1052_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3161 _1052_/a_891_413# _1052_/a_27_47# _1052_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3162 _1052_/a_592_47# _1052_/a_193_47# _1052_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3163 VPWR _1052_/a_1059_315# _1052_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3164 _1052_/a_1017_47# _1052_/a_27_47# _1052_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3165 _1052_/a_193_47# _1052_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3166 _1052_/a_466_413# _1052_/a_27_47# _1052_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3167 VGND _1052_/a_891_413# _1052_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3168 _1052_/a_381_47# _0150_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3169 VGND net138 _1052_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3170 VGND _0218_ _0836_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X3171 _0836_/a_68_297# net248 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3172 _0442_ _0836_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3173 VPWR _0218_ _0836_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X3174 _0442_ _0836_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X3175 _0836_/a_150_297# net248 _0836_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3176 VPWR _0305_ _0767_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X3177 _0387_ _0767_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X3178 VGND _0305_ _0767_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X3179 _0767_/a_59_75# _0294_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3180 _0387_ _0767_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X3181 _0767_/a_145_75# _0294_ _0767_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X3182 _0698_/a_199_47# _0317_ _0330_ VGND sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.182 ps=1.86 w=0.65 l=0.15
X3183 _0698_/a_113_297# _0319_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.545 pd=5.09 as=0 ps=0 w=1 l=0.15
X3184 _0330_ _0316_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3185 VPWR _0317_ _0698_/a_113_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3186 _0698_/a_113_297# _0316_ _0330_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X3187 VGND _0319_ _0698_/a_199_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3188 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3189 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3190 _0253_ _0621_/a_35_297# _0621_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.53 ps=5.06 w=1 l=0.15
X3191 _0253_ net64 _0621_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.5005 pd=2.84 as=0.1755 ps=1.84 w=0.65 l=0.15
X3192 _0621_/a_35_297# net64 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X3193 _0621_/a_117_297# net64 _0621_/a_35_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.26 ps=2.52 w=1 l=0.15
X3194 VPWR net64 _0621_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3195 VGND acc0.A\[6\] _0621_/a_35_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3196 VGND _0621_/a_35_297# _0253_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3197 _0621_/a_285_297# acc0.A\[6\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3198 VPWR acc0.A\[6\] _0621_/a_117_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3199 _0621_/a_285_47# acc0.A\[6\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3200 VGND comp0.B\[6\] _0552_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X3201 _0552_/a_68_297# _0176_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3202 _0209_ _0552_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3203 VPWR comp0.B\[6\] _0552_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X3204 _0209_ _0552_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X3205 _0552_/a_150_297# _0176_ _0552_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3206 comp0.B\[3\] _1035_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3207 _1035_/a_891_413# _1035_/a_193_47# _1035_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3208 _1035_/a_561_413# _1035_/a_27_47# _1035_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3209 VPWR net121 _1035_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3210 comp0.B\[3\] _1035_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3211 _1035_/a_381_47# _0133_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3212 VGND _1035_/a_634_159# _1035_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3213 VPWR _1035_/a_891_413# _1035_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3214 _1035_/a_466_413# _1035_/a_193_47# _1035_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3215 VPWR _1035_/a_634_159# _1035_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3216 _1035_/a_634_159# _1035_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3217 _1035_/a_634_159# _1035_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3218 _1035_/a_975_413# _1035_/a_193_47# _1035_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3219 VGND _1035_/a_1059_315# _1035_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3220 _1035_/a_193_47# _1035_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3221 _1035_/a_891_413# _1035_/a_27_47# _1035_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3222 _1035_/a_592_47# _1035_/a_193_47# _1035_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3223 VPWR _1035_/a_1059_315# _1035_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3224 _1035_/a_1017_47# _1035_/a_27_47# _1035_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3225 _1035_/a_193_47# _1035_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3226 _1035_/a_466_413# _1035_/a_27_47# _1035_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3227 VGND _1035_/a_891_413# _1035_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3228 _1035_/a_381_47# _0133_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3229 VGND net121 _1035_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3230 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3231 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3232 _0819_/a_81_21# _0346_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X3233 _0819_/a_299_297# _0346_ _0819_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X3234 VPWR _0819_/a_81_21# _0428_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X3235 VPWR _0401_ _0819_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3236 VGND _0819_/a_81_21# _0428_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3237 VGND _0427_ _0819_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X3238 _0819_/a_299_297# _0427_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3239 _0819_/a_384_47# _0401_ _0819_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3240 net92 clknet_1_0__leaf__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X3241 VGND clknet_1_0__leaf__0460_ net92 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X3242 net92 clknet_1_0__leaf__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3243 VPWR clknet_1_0__leaf__0460_ net92 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3244 VPWR _0226_ _0236_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3245 _0236_ _0226_ _0604_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X3246 _0604_/a_113_47# _0235_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3247 _0236_ _0235_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3248 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3249 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3250 VGND comp0.B\[14\] _0535_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X3251 _0535_/a_68_297# _0176_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3252 _0200_ _0535_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3253 VPWR comp0.B\[14\] _0535_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X3254 _0200_ _0535_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X3255 _0535_/a_150_297# _0176_ _0535_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3256 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3257 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3258 acc0.A\[18\] _1018_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3259 _1018_/a_891_413# _1018_/a_193_47# _1018_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3260 _1018_/a_561_413# _1018_/a_27_47# _1018_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3261 VPWR net104 _1018_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3262 acc0.A\[18\] _1018_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3263 _1018_/a_381_47# _0116_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3264 VGND _1018_/a_634_159# _1018_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3265 VPWR _1018_/a_891_413# _1018_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3266 _1018_/a_466_413# _1018_/a_193_47# _1018_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3267 VPWR _1018_/a_634_159# _1018_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3268 _1018_/a_634_159# _1018_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3269 _1018_/a_634_159# _1018_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3270 _1018_/a_975_413# _1018_/a_193_47# _1018_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3271 VGND _1018_/a_1059_315# _1018_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3272 _1018_/a_193_47# _1018_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3273 _1018_/a_891_413# _1018_/a_27_47# _1018_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3274 _1018_/a_592_47# _1018_/a_193_47# _1018_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3275 VPWR _1018_/a_1059_315# _1018_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3276 _1018_/a_1017_47# _1018_/a_27_47# _1018_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3277 _1018_/a_193_47# _1018_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3278 _1018_/a_466_413# _1018_/a_27_47# _1018_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3279 VGND _1018_/a_891_413# _1018_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3280 _1018_/a_381_47# _0116_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3281 VGND net104 _1018_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3282 VPWR clknet_0__0464_ clkbuf_1_1__f__0464_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X3283 VPWR clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X3284 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3285 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3286 VPWR clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3287 VPWR clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3288 clkbuf_1_1__f__0464_/a_110_47# clknet_0__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3289 clkbuf_1_1__f__0464_/a_110_47# clknet_0__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X3290 VGND clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X3291 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3292 VGND clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3293 clkbuf_1_1__f__0464_/a_110_47# clknet_0__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3294 VGND clknet_0__0464_ clkbuf_1_1__f__0464_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3295 VGND clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3296 VPWR clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3297 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3298 VGND clknet_0__0464_ clkbuf_1_1__f__0464_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3299 VGND clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3300 VPWR clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3301 VGND clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3302 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3303 clkbuf_1_1__f__0464_/a_110_47# clknet_0__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3304 VPWR clknet_0__0464_ clkbuf_1_1__f__0464_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3305 VPWR clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3306 VPWR clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3307 VGND clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3308 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3309 VGND clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3310 VGND clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3311 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3312 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3313 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3314 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3315 VPWR clkbuf_1_1__f__0464_/a_110_47# clknet_1_1__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3316 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3317 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3318 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3319 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3320 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3321 clknet_1_1__leaf__0464_ clkbuf_1_1__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3322 VPWR net15 _0518_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X3323 _0518_/a_27_297# _0186_ _0518_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X3324 VGND net15 _0518_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X3325 _0191_ _0518_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3326 _0518_/a_27_297# _0186_ _0518_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X3327 _0518_/a_109_297# _0180_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3328 _0518_/a_373_47# _0180_ _0518_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3329 _0191_ _0518_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3330 _0518_/a_109_297# acc0.A\[8\] _0518_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3331 _0518_/a_109_47# acc0.A\[8\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3332 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3333 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3334 net43 _0998_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3335 _0998_/a_891_413# _0998_/a_193_47# _0998_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3336 _0998_/a_561_413# _0998_/a_27_47# _0998_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3337 VPWR net84 _0998_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3338 net43 _0998_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3339 _0998_/a_381_47# _0096_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3340 VGND _0998_/a_634_159# _0998_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3341 VPWR _0998_/a_891_413# _0998_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3342 _0998_/a_466_413# _0998_/a_193_47# _0998_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3343 VPWR _0998_/a_634_159# _0998_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3344 _0998_/a_634_159# _0998_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3345 _0998_/a_634_159# _0998_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3346 _0998_/a_975_413# _0998_/a_193_47# _0998_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3347 VGND _0998_/a_1059_315# _0998_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3348 _0998_/a_193_47# _0998_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3349 _0998_/a_891_413# _0998_/a_27_47# _0998_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3350 _0998_/a_592_47# _0998_/a_193_47# _0998_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3351 VPWR _0998_/a_1059_315# _0998_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3352 _0998_/a_1017_47# _0998_/a_27_47# _0998_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3353 _0998_/a_193_47# _0998_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3354 _0998_/a_466_413# _0998_/a_27_47# _0998_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3355 VGND _0998_/a_891_413# _0998_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3356 _0998_/a_381_47# _0096_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3357 VGND net84 _0998_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3358 _0454_ _0852_/a_35_297# _0852_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.53 ps=5.06 w=1 l=0.15
X3359 _0454_ _0453_ _0852_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.5005 pd=2.84 as=0.1755 ps=1.84 w=0.65 l=0.15
X3360 _0852_/a_35_297# _0453_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X3361 _0852_/a_117_297# _0453_ _0852_/a_35_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.26 ps=2.52 w=1 l=0.15
X3362 VPWR _0453_ _0852_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3363 VGND _0264_ _0852_/a_35_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3364 VGND _0852_/a_35_297# _0454_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3365 _0852_/a_285_297# _0264_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3366 VPWR _0264_ _0852_/a_117_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3367 _0852_/a_285_47# _0264_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3368 VGND _0347_ _0783_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X3369 _0783_/a_510_47# _0398_ _0783_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X3370 _0783_/a_79_21# _0399_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X3371 VPWR _0398_ _0783_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3372 _0783_/a_79_21# _0397_ _0783_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X3373 _0783_/a_297_297# _0347_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3374 _0783_/a_79_21# _0399_ _0783_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X3375 VPWR _0783_/a_79_21# _0096_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X3376 VGND _0783_/a_79_21# _0096_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3377 _0783_/a_215_47# _0397_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3378 VPWR input2/a_75_212# net2 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X3379 input2/a_75_212# A[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X3380 input2/a_75_212# A[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3381 VGND input2/a_75_212# net2 VGND sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X3382 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X3383 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X3384 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X3385 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X3386 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3387 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3388 acc0.A\[5\] _1051_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3389 _1051_/a_891_413# _1051_/a_193_47# _1051_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3390 _1051_/a_561_413# _1051_/a_27_47# _1051_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3391 VPWR net137 _1051_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3392 acc0.A\[5\] _1051_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3393 _1051_/a_381_47# _0149_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3394 VGND _1051_/a_634_159# _1051_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3395 VPWR _1051_/a_891_413# _1051_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3396 _1051_/a_466_413# _1051_/a_193_47# _1051_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3397 VPWR _1051_/a_634_159# _1051_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3398 _1051_/a_634_159# _1051_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3399 _1051_/a_634_159# _1051_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3400 _1051_/a_975_413# _1051_/a_193_47# _1051_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3401 VGND _1051_/a_1059_315# _1051_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3402 _1051_/a_193_47# _1051_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3403 _1051_/a_891_413# _1051_/a_27_47# _1051_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3404 _1051_/a_592_47# _1051_/a_193_47# _1051_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3405 VPWR _1051_/a_1059_315# _1051_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3406 _1051_/a_1017_47# _1051_/a_27_47# _1051_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3407 _1051_/a_193_47# _1051_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3408 _1051_/a_466_413# _1051_/a_27_47# _1051_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3409 VGND _1051_/a_891_413# _1051_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3410 _1051_/a_381_47# _0149_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3411 VGND net137 _1051_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3412 _0835_/a_78_199# _0432_ _0835_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3413 VPWR _0257_ _0835_/a_493_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X3414 _0835_/a_493_297# _0255_ _0835_/a_78_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.235 ps=1.47 w=1 l=0.15
X3415 VPWR _0835_/a_78_199# _0441_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3725 pd=1.745 as=0.28 ps=2.56 w=1 l=0.15
X3416 VGND _0255_ _0835_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.11375 ps=1 w=0.65 l=0.15
X3417 _0835_/a_78_199# _0256_ _0835_/a_292_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.235 pd=1.47 as=0.1175 ps=1.235 w=1 l=0.15
X3418 _0835_/a_215_47# _0257_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3419 _0835_/a_215_47# _0256_ _0835_/a_78_199# VGND sky130_fd_pr__nfet_01v8 ad=0.11375 pd=1 as=0.08775 ps=0.92 w=0.65 l=0.15
X3420 _0835_/a_292_297# _0432_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1175 pd=1.235 as=0.3725 ps=1.745 w=1 l=0.15
X3421 VGND _0835_/a_78_199# _0441_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X3422 VPWR _0244_ _0766_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X3423 VGND _0244_ _0386_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X3424 _0766_/a_109_297# _0245_ _0386_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X3425 _0386_ _0245_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3426 VPWR _0697_/a_80_21# _0329_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X3427 _0697_/a_80_21# _0322_ _0697_/a_472_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.31 ps=2.62 w=1 l=0.15
X3428 VPWR _0313_ _0697_/a_217_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.545 ps=5.09 w=1 l=0.15
X3429 VGND _0328_ _0697_/a_80_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.35425 ps=3.69 w=0.65 l=0.15
X3430 VGND _0697_/a_80_21# _0329_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.17225 ps=1.83 w=0.65 l=0.15
X3431 _0697_/a_300_47# _0313_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X3432 _0697_/a_217_297# _0324_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3433 _0697_/a_80_21# _0324_ _0697_/a_300_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3434 _0697_/a_472_297# _0328_ _0697_/a_217_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3435 _0697_/a_80_21# _0322_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3436 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3437 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3438 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3439 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3440 VPWR acc0.A\[7\] _0252_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3441 _0252_ acc0.A\[7\] _0620_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X3442 _0620_/a_113_47# net65 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3443 _0252_ net65 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3444 VPWR _0551_/a_27_47# _0208_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3445 _0208_ _0551_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3446 VPWR _0171_ _0551_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3447 _0208_ _0551_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X3448 VGND _0551_/a_27_47# _0208_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3449 VGND _0171_ _0551_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3450 comp0.B\[2\] _1034_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3451 _1034_/a_891_413# _1034_/a_193_47# _1034_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3452 _1034_/a_561_413# _1034_/a_27_47# _1034_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3453 VPWR net120 _1034_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3454 comp0.B\[2\] _1034_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3455 _1034_/a_381_47# net186 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3456 VGND _1034_/a_634_159# _1034_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3457 VPWR _1034_/a_891_413# _1034_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3458 _1034_/a_466_413# _1034_/a_193_47# _1034_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3459 VPWR _1034_/a_634_159# _1034_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3460 _1034_/a_634_159# _1034_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3461 _1034_/a_634_159# _1034_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3462 _1034_/a_975_413# _1034_/a_193_47# _1034_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3463 VGND _1034_/a_1059_315# _1034_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3464 _1034_/a_193_47# _1034_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3465 _1034_/a_891_413# _1034_/a_27_47# _1034_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3466 _1034_/a_592_47# _1034_/a_193_47# _1034_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3467 VPWR _1034_/a_1059_315# _1034_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3468 _1034_/a_1017_47# _1034_/a_27_47# _1034_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3469 _1034_/a_193_47# _1034_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3470 _1034_/a_466_413# _1034_/a_27_47# _1034_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3471 VGND _1034_/a_891_413# _1034_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3472 _1034_/a_381_47# net186 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3473 VGND net120 _1034_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3474 VPWR _0275_ _0427_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.53 ps=5.06 w=1 l=0.15
X3475 _0427_ _0259_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3476 _0818_/a_193_47# _0275_ _0818_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.1755 ps=1.84 w=0.65 l=0.15
X3477 _0427_ _0259_ _0818_/a_193_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3478 _0427_ _0292_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3479 _0818_/a_109_47# _0292_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3480 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3481 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3482 _0749_/a_81_21# _0236_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X3483 _0749_/a_299_297# _0236_ _0749_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X3484 VPWR _0749_/a_81_21# _0373_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X3485 VPWR _0248_ _0749_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3486 VGND _0749_/a_81_21# _0373_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3487 VGND _0372_ _0749_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X3488 _0749_/a_299_297# _0372_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3489 _0749_/a_384_47# _0248_ _0749_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3490 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3491 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3492 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3493 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3494 _0534_/a_81_21# _0199_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X3495 _0534_/a_299_297# _0199_ _0534_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X3496 VPWR _0534_/a_81_21# _0145_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X3497 VPWR net149 _0534_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3498 VGND _0534_/a_81_21# _0145_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3499 VGND _0195_ _0534_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X3500 _0534_/a_299_297# _0195_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3501 _0534_/a_384_47# net149 _0534_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3502 VGND acc0.A\[20\] _0603_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X3503 _0603_/a_68_297# net48 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3504 _0235_ _0603_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3505 VPWR acc0.A\[20\] _0603_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X3506 _0235_ _0603_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X3507 _0603_/a_150_297# net48 _0603_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3508 acc0.A\[17\] _1017_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3509 _1017_/a_891_413# _1017_/a_193_47# _1017_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3510 _1017_/a_561_413# _1017_/a_27_47# _1017_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3511 VPWR net103 _1017_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3512 acc0.A\[17\] _1017_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3513 _1017_/a_381_47# _0115_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3514 VGND _1017_/a_634_159# _1017_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3515 VPWR _1017_/a_891_413# _1017_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3516 _1017_/a_466_413# _1017_/a_193_47# _1017_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3517 VPWR _1017_/a_634_159# _1017_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3518 _1017_/a_634_159# _1017_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3519 _1017_/a_634_159# _1017_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3520 _1017_/a_975_413# _1017_/a_193_47# _1017_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3521 VGND _1017_/a_1059_315# _1017_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3522 _1017_/a_193_47# _1017_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3523 _1017_/a_891_413# _1017_/a_27_47# _1017_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3524 _1017_/a_592_47# _1017_/a_193_47# _1017_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3525 VPWR _1017_/a_1059_315# _1017_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3526 _1017_/a_1017_47# _1017_/a_27_47# _1017_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3527 _1017_/a_193_47# _1017_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3528 _1017_/a_466_413# _1017_/a_27_47# _1017_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3529 VGND _1017_/a_891_413# _1017_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3530 _1017_/a_381_47# _0115_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3531 VGND net103 _1017_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3532 VPWR clknet_0__0463_ clkbuf_1_1__f__0463_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X3533 VPWR clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X3534 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3535 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3536 VPWR clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3537 VPWR clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3538 clkbuf_1_1__f__0463_/a_110_47# clknet_0__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3539 clkbuf_1_1__f__0463_/a_110_47# clknet_0__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X3540 VGND clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X3541 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3542 VGND clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3543 clkbuf_1_1__f__0463_/a_110_47# clknet_0__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3544 VGND clknet_0__0463_ clkbuf_1_1__f__0463_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3545 VGND clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3546 VPWR clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3547 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3548 VGND clknet_0__0463_ clkbuf_1_1__f__0463_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3549 VGND clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3550 VPWR clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3551 VGND clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3552 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3553 clkbuf_1_1__f__0463_/a_110_47# clknet_0__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3554 VPWR clknet_0__0463_ clkbuf_1_1__f__0463_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3555 VPWR clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3556 VPWR clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3557 VGND clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3558 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3559 VGND clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3560 VGND clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3561 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3562 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3563 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3564 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3565 VPWR clkbuf_1_1__f__0463_/a_110_47# clknet_1_1__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3566 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3567 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3568 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3569 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3570 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3571 clknet_1_1__leaf__0463_ clkbuf_1_1__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3572 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3573 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3574 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3575 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3576 _0517_/a_81_21# _0190_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X3577 _0517_/a_299_297# _0190_ _0517_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X3578 VPWR _0517_/a_81_21# _0153_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X3579 VPWR net178 _0517_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3580 VGND _0517_/a_81_21# _0153_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3581 VGND _0179_ _0517_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X3582 _0517_/a_299_297# _0179_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3583 _0517_/a_384_47# net178 _0517_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3584 net130 clknet_1_1__leaf__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X3585 VGND clknet_1_1__leaf__0464_ net130 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X3586 net130 clknet_1_1__leaf__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3587 VPWR clknet_1_1__leaf__0464_ net130 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3588 net144 clknet_1_1__leaf__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X3589 VGND clknet_1_1__leaf__0465_ net144 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X3590 net144 clknet_1_1__leaf__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3591 VPWR clknet_1_1__leaf__0465_ net144 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3592 net42 _0997_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3593 _0997_/a_891_413# _0997_/a_193_47# _0997_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3594 _0997_/a_561_413# _0997_/a_27_47# _0997_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3595 VPWR net83 _0997_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3596 net42 _0997_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3597 _0997_/a_381_47# _0095_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3598 VGND _0997_/a_634_159# _0997_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3599 VPWR _0997_/a_891_413# _0997_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3600 _0997_/a_466_413# _0997_/a_193_47# _0997_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3601 VPWR _0997_/a_634_159# _0997_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3602 _0997_/a_634_159# _0997_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3603 _0997_/a_634_159# _0997_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3604 _0997_/a_975_413# _0997_/a_193_47# _0997_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3605 VGND _0997_/a_1059_315# _0997_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3606 _0997_/a_193_47# _0997_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3607 _0997_/a_891_413# _0997_/a_27_47# _0997_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3608 _0997_/a_592_47# _0997_/a_193_47# _0997_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3609 VPWR _0997_/a_1059_315# _0997_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3610 _0997_/a_1017_47# _0997_/a_27_47# _0997_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3611 _0997_/a_193_47# _0997_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3612 _0997_/a_466_413# _0997_/a_27_47# _0997_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3613 VGND _0997_/a_891_413# _0997_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3614 _0997_/a_381_47# _0095_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3615 VGND net83 _0997_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3616 VPWR _0465_ clkbuf_0__0465_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X3617 VPWR clkbuf_0__0465_/a_110_47# clknet_0__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X3618 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3619 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3620 VPWR clkbuf_0__0465_/a_110_47# clknet_0__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3621 VPWR clkbuf_0__0465_/a_110_47# clknet_0__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3622 clkbuf_0__0465_/a_110_47# _0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3623 clkbuf_0__0465_/a_110_47# _0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X3624 VGND clkbuf_0__0465_/a_110_47# clknet_0__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X3625 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3626 VGND clkbuf_0__0465_/a_110_47# clknet_0__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3627 clkbuf_0__0465_/a_110_47# _0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3628 VGND _0465_ clkbuf_0__0465_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3629 VGND clkbuf_0__0465_/a_110_47# clknet_0__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3630 VPWR clkbuf_0__0465_/a_110_47# clknet_0__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3631 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3632 VGND _0465_ clkbuf_0__0465_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3633 VGND clkbuf_0__0465_/a_110_47# clknet_0__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3634 VPWR clkbuf_0__0465_/a_110_47# clknet_0__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3635 VGND clkbuf_0__0465_/a_110_47# clknet_0__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3636 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3637 clkbuf_0__0465_/a_110_47# _0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3638 VPWR _0465_ clkbuf_0__0465_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3639 VPWR clkbuf_0__0465_/a_110_47# clknet_0__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3640 VPWR clkbuf_0__0465_/a_110_47# clknet_0__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3641 VGND clkbuf_0__0465_/a_110_47# clknet_0__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3642 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3643 VGND clkbuf_0__0465_/a_110_47# clknet_0__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3644 VGND clkbuf_0__0465_/a_110_47# clknet_0__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3645 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3646 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3647 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3648 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3649 VPWR clkbuf_0__0465_/a_110_47# clknet_0__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3650 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3651 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3652 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3653 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3654 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3655 clknet_0__0465_ clkbuf_0__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3656 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3657 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3658 VPWR _0266_ _0453_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3659 _0453_ _0266_ _0851_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X3660 _0851_/a_113_47# _0452_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3661 _0453_ _0452_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3662 VPWR _0208_ _0782_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X3663 VGND _0782_/a_27_47# _0399_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X3664 VGND _0782_/a_27_47# _0399_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3665 _0399_ _0782_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X3666 _0399_ _0782_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3667 VGND _0208_ _0782_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X3668 VPWR _0782_/a_27_47# _0399_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3669 _0399_ _0782_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3670 _0399_ _0782_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3671 VPWR _0782_/a_27_47# _0399_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3672 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3673 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3674 net111 clknet_1_0__leaf__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X3675 VGND clknet_1_0__leaf__0462_ net111 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X3676 net111 clknet_1_0__leaf__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3677 VPWR clknet_1_0__leaf__0462_ net111 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3678 net125 clknet_1_0__leaf__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X3679 VGND clknet_1_0__leaf__0463_ net125 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X3680 net125 clknet_1_0__leaf__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3681 VPWR clknet_1_0__leaf__0463_ net125 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3682 VPWR input3/a_75_212# net3 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X3683 input3/a_75_212# A[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X3684 input3/a_75_212# A[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X3685 VGND input3/a_75_212# net3 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X3686 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3687 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3688 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3689 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3690 acc0.A\[4\] _1050_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3691 _1050_/a_891_413# _1050_/a_193_47# _1050_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3692 _1050_/a_561_413# _1050_/a_27_47# _1050_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3693 VPWR net136 _1050_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3694 acc0.A\[4\] _1050_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3695 _1050_/a_381_47# _0148_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3696 VGND _1050_/a_634_159# _1050_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3697 VPWR _1050_/a_891_413# _1050_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3698 _1050_/a_466_413# _1050_/a_193_47# _1050_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3699 VPWR _1050_/a_634_159# _1050_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3700 _1050_/a_634_159# _1050_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3701 _1050_/a_634_159# _1050_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3702 _1050_/a_975_413# _1050_/a_193_47# _1050_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3703 VGND _1050_/a_1059_315# _1050_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3704 _1050_/a_193_47# _1050_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3705 _1050_/a_891_413# _1050_/a_27_47# _1050_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3706 _1050_/a_592_47# _1050_/a_193_47# _1050_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3707 VPWR _1050_/a_1059_315# _1050_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3708 _1050_/a_1017_47# _1050_/a_27_47# _1050_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3709 _1050_/a_193_47# _1050_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3710 _1050_/a_466_413# _1050_/a_27_47# _1050_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3711 VGND _1050_/a_891_413# _1050_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3712 _1050_/a_381_47# _0148_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3713 VGND net136 _1050_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3714 VPWR _0255_ _0834_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X3715 VGND _0255_ _0440_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X3716 _0834_/a_109_297# _0433_ _0440_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X3717 _0440_ _0433_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3718 VPWR acc0.A\[25\] _0696_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X3719 VGND acc0.A\[25\] _0328_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X3720 _0696_/a_109_297# net53 _0328_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X3721 _0328_ net53 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3722 VGND _0369_ _0765_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X3723 _0765_/a_510_47# _0385_ _0765_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X3724 _0765_/a_79_21# _0352_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X3725 VPWR _0385_ _0765_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3726 _0765_/a_79_21# net220 _0765_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X3727 _0765_/a_297_297# _0369_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3728 _0765_/a_79_21# _0352_ _0765_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X3729 VPWR _0765_/a_79_21# _0100_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X3730 VGND _0765_/a_79_21# _0100_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3731 _0765_/a_215_47# net220 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3732 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3733 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3734 net106 clknet_1_0__leaf__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X3735 VGND clknet_1_0__leaf__0461_ net106 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X3736 net106 clknet_1_0__leaf__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3737 VPWR clknet_1_0__leaf__0461_ net106 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3738 _0550_/a_240_47# net30 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X3739 _0137_ _0550_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X3740 VGND _0172_ _0550_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3741 _0550_/a_51_297# net180 _0550_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X3742 _0550_/a_149_47# _0207_ _0550_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X3743 _0550_/a_240_47# _0174_ _0550_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3744 VPWR _0172_ _0550_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X3745 _0137_ _0550_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X3746 _0550_/a_149_47# net180 _0550_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3747 _0550_/a_245_297# _0174_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3748 VPWR _0207_ _0550_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3749 _0550_/a_512_297# net30 _0550_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3750 comp0.B\[1\] _1033_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3751 _1033_/a_891_413# _1033_/a_193_47# _1033_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3752 _1033_/a_561_413# _1033_/a_27_47# _1033_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3753 VPWR net119 _1033_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3754 comp0.B\[1\] _1033_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3755 _1033_/a_381_47# _0131_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3756 VGND _1033_/a_634_159# _1033_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3757 VPWR _1033_/a_891_413# _1033_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3758 _1033_/a_466_413# _1033_/a_193_47# _1033_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3759 VPWR _1033_/a_634_159# _1033_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3760 _1033_/a_634_159# _1033_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3761 _1033_/a_634_159# _1033_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3762 _1033_/a_975_413# _1033_/a_193_47# _1033_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3763 VGND _1033_/a_1059_315# _1033_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3764 _1033_/a_193_47# _1033_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3765 _1033_/a_891_413# _1033_/a_27_47# _1033_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3766 _1033_/a_592_47# _1033_/a_193_47# _1033_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3767 VPWR _1033_/a_1059_315# _1033_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3768 _1033_/a_1017_47# _1033_/a_27_47# _1033_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3769 _1033_/a_193_47# _1033_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3770 _1033_/a_466_413# _1033_/a_27_47# _1033_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3771 VGND _1033_/a_891_413# _1033_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3772 _1033_/a_381_47# _0131_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3773 VGND net119 _1033_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3774 _0817_/a_585_47# _0426_ _0817_/a_266_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.72 as=0.47125 ps=4.05 w=0.65 l=0.15
X3775 VGND _0424_ _0817_/a_266_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3776 VPWR _0817_/a_81_21# _0089_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X3777 _0817_/a_81_21# _0345_ _0817_/a_585_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3778 VGND _0817_/a_81_21# _0089_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3779 _0817_/a_266_297# _0346_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0 ps=0 w=1 l=0.15
X3780 _0817_/a_368_297# _0424_ _0817_/a_266_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.42 pd=2.84 as=0 ps=0 w=1 l=0.15
X3781 _0817_/a_266_47# _0425_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3782 _0817_/a_266_47# _0346_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3783 _0817_/a_81_21# _0425_ _0817_/a_368_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.535 pd=5.07 as=0 ps=0 w=1 l=0.15
X3784 _0817_/a_81_21# _0345_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3785 VPWR _0426_ _0817_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3786 _0748_/a_81_21# _0311_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X3787 _0748_/a_299_297# _0311_ _0748_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X3788 VPWR _0748_/a_81_21# _0372_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X3789 VPWR _0294_ _0748_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3790 VGND _0748_/a_81_21# _0372_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3791 VGND _0305_ _0748_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X3792 _0748_/a_299_297# _0305_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3793 _0748_/a_384_47# _0294_ _0748_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3794 VGND _0246_ _0679_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X3795 _0679_/a_68_297# _0310_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3796 _0311_ _0679_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3797 VPWR _0246_ _0679_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X3798 _0311_ _0679_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X3799 _0679_/a_150_297# _0310_ _0679_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3800 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3801 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3802 VPWR _0233_ _0234_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3803 _0234_ _0233_ _0602_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X3804 _0602_/a_113_47# _0231_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3805 _0234_ _0231_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3806 VPWR net8 _0533_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X3807 _0533_/a_27_297# _0182_ _0533_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X3808 VGND net8 _0533_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X3809 _0199_ _0533_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3810 _0533_/a_27_297# _0182_ _0533_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X3811 _0533_/a_109_297# _0180_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3812 _0533_/a_373_47# _0180_ _0533_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3813 _0199_ _0533_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3814 _0533_/a_109_297# acc0.A\[1\] _0533_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3815 _0533_/a_109_47# acc0.A\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3816 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X3817 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X3818 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3819 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3820 acc0.A\[16\] _1016_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3821 _1016_/a_891_413# _1016_/a_193_47# _1016_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3822 _1016_/a_561_413# _1016_/a_27_47# _1016_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3823 VPWR net102 _1016_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3824 acc0.A\[16\] _1016_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3825 _1016_/a_381_47# net166 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3826 VGND _1016_/a_634_159# _1016_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3827 VPWR _1016_/a_891_413# _1016_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3828 _1016_/a_466_413# _1016_/a_193_47# _1016_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3829 VPWR _1016_/a_634_159# _1016_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3830 _1016_/a_634_159# _1016_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3831 _1016_/a_634_159# _1016_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3832 _1016_/a_975_413# _1016_/a_193_47# _1016_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3833 VGND _1016_/a_1059_315# _1016_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3834 _1016_/a_193_47# _1016_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3835 _1016_/a_891_413# _1016_/a_27_47# _1016_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3836 _1016_/a_592_47# _1016_/a_193_47# _1016_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3837 VPWR _1016_/a_1059_315# _1016_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3838 _1016_/a_1017_47# _1016_/a_27_47# _1016_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3839 _1016_/a_193_47# _1016_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3840 _1016_/a_466_413# _1016_/a_27_47# _1016_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3841 VGND _1016_/a_891_413# _1016_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3842 _1016_/a_381_47# net166 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3843 VGND net102 _1016_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3844 VPWR clknet_0__0462_ clkbuf_1_1__f__0462_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X3845 VPWR clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X3846 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3847 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3848 VPWR clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3849 VPWR clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3850 clkbuf_1_1__f__0462_/a_110_47# clknet_0__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3851 clkbuf_1_1__f__0462_/a_110_47# clknet_0__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X3852 VGND clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X3853 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3854 VGND clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3855 clkbuf_1_1__f__0462_/a_110_47# clknet_0__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3856 VGND clknet_0__0462_ clkbuf_1_1__f__0462_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3857 VGND clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3858 VPWR clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3859 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3860 VGND clknet_0__0462_ clkbuf_1_1__f__0462_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3861 VGND clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3862 VPWR clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3863 VGND clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3864 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3865 clkbuf_1_1__f__0462_/a_110_47# clknet_0__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3866 VPWR clknet_0__0462_ clkbuf_1_1__f__0462_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3867 VPWR clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3868 VPWR clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3869 VGND clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3870 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3871 VGND clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3872 VGND clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3873 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3874 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3875 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3876 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3877 VPWR clkbuf_1_1__f__0462_/a_110_47# clknet_1_1__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3878 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3879 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3880 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3881 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3882 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3883 clknet_1_1__leaf__0462_ clkbuf_1_1__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3884 net97 clknet_1_1__leaf__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X3885 VGND clknet_1_1__leaf__0460_ net97 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X3886 net97 clknet_1_1__leaf__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3887 VPWR clknet_1_1__leaf__0460_ net97 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3888 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3889 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3890 VPWR net16 _0516_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X3891 _0516_/a_27_297# _0186_ _0516_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X3892 VGND net16 _0516_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X3893 _0190_ _0516_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3894 _0516_/a_27_297# _0186_ _0516_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X3895 _0516_/a_109_297# _0181_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3896 _0516_/a_373_47# _0181_ _0516_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3897 _0190_ _0516_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3898 _0516_/a_109_297# acc0.A\[9\] _0516_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3899 _0516_/a_109_47# acc0.A\[9\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X3900 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X3901 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X3902 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X3903 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X3904 net41 _0996_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3905 _0996_/a_891_413# _0996_/a_193_47# _0996_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X3906 _0996_/a_561_413# _0996_/a_27_47# _0996_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X3907 VPWR net82 _0996_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X3908 net41 _0996_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X3909 _0996_/a_381_47# _0094_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X3910 VGND _0996_/a_634_159# _0996_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X3911 VPWR _0996_/a_891_413# _0996_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X3912 _0996_/a_466_413# _0996_/a_193_47# _0996_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3913 VPWR _0996_/a_634_159# _0996_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3914 _0996_/a_634_159# _0996_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X3915 _0996_/a_634_159# _0996_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X3916 _0996_/a_975_413# _0996_/a_193_47# _0996_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X3917 VGND _0996_/a_1059_315# _0996_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X3918 _0996_/a_193_47# _0996_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X3919 _0996_/a_891_413# _0996_/a_27_47# _0996_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3920 _0996_/a_592_47# _0996_/a_193_47# _0996_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X3921 VPWR _0996_/a_1059_315# _0996_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3922 _0996_/a_1017_47# _0996_/a_27_47# _0996_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X3923 _0996_/a_193_47# _0996_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X3924 _0996_/a_466_413# _0996_/a_27_47# _0996_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X3925 VGND _0996_/a_891_413# _0996_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X3926 _0996_/a_381_47# _0094_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3927 VGND net82 _0996_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3928 VPWR _0464_ clkbuf_0__0464_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X3929 VPWR clkbuf_0__0464_/a_110_47# clknet_0__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X3930 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3931 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3932 VPWR clkbuf_0__0464_/a_110_47# clknet_0__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3933 VPWR clkbuf_0__0464_/a_110_47# clknet_0__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3934 clkbuf_0__0464_/a_110_47# _0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3935 clkbuf_0__0464_/a_110_47# _0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X3936 VGND clkbuf_0__0464_/a_110_47# clknet_0__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X3937 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3938 VGND clkbuf_0__0464_/a_110_47# clknet_0__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3939 clkbuf_0__0464_/a_110_47# _0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3940 VGND _0464_ clkbuf_0__0464_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3941 VGND clkbuf_0__0464_/a_110_47# clknet_0__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3942 VPWR clkbuf_0__0464_/a_110_47# clknet_0__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3943 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3944 VGND _0464_ clkbuf_0__0464_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3945 VGND clkbuf_0__0464_/a_110_47# clknet_0__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3946 VPWR clkbuf_0__0464_/a_110_47# clknet_0__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3947 VGND clkbuf_0__0464_/a_110_47# clknet_0__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3948 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3949 clkbuf_0__0464_/a_110_47# _0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3950 VPWR _0464_ clkbuf_0__0464_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3951 VPWR clkbuf_0__0464_/a_110_47# clknet_0__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3952 VPWR clkbuf_0__0464_/a_110_47# clknet_0__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3953 VGND clkbuf_0__0464_/a_110_47# clknet_0__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3954 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3955 VGND clkbuf_0__0464_/a_110_47# clknet_0__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3956 VGND clkbuf_0__0464_/a_110_47# clknet_0__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3957 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3958 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3959 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3960 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3961 VPWR clkbuf_0__0464_/a_110_47# clknet_0__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3962 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X3963 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3964 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3965 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3966 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3967 clknet_0__0464_ clkbuf_0__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3968 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3969 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3970 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3971 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3972 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3973 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3974 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3975 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3976 VGND acc0.A\[1\] _0850_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X3977 _0850_/a_68_297# net47 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3978 _0452_ _0850_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3979 VPWR acc0.A\[1\] _0850_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X3980 _0452_ _0850_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X3981 _0850_/a_150_297# net47 _0850_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3982 VGND _0218_ _0781_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X3983 _0781_/a_68_297# net43 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X3984 _0398_ _0781_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X3985 VPWR _0218_ _0781_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X3986 _0398_ _0781_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X3987 _0781_/a_150_297# net43 _0781_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X3988 VPWR input4/a_75_212# net4 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X3989 input4/a_75_212# A[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X3990 input4/a_75_212# A[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X3991 VGND input4/a_75_212# net4 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X3992 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X3993 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X3994 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X3995 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X3996 VPWR _0466_ _0979_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X3997 _0979_/a_27_297# _0480_ _0979_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X3998 VGND _0466_ _0979_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X3999 _0169_ _0979_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4000 _0979_/a_27_297# _0480_ _0979_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X4001 _0979_/a_109_297# net164 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4002 _0979_/a_373_47# net164 _0979_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4003 _0169_ _0979_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4004 _0979_/a_109_297# _0488_ _0979_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4005 _0979_/a_109_47# _0488_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4006 VPWR clknet_1_0__leaf__0457_ _0902_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X4007 _0462_ _0902_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X4008 _0462_ _0902_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X4009 VGND clknet_1_0__leaf__0457_ _0902_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X4010 VGND _0369_ _0833_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X4011 _0833_/a_510_47# _0439_ _0833_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X4012 _0833_/a_79_21# _0399_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X4013 VPWR _0439_ _0833_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4014 _0833_/a_79_21# net235 _0833_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X4015 _0833_/a_297_297# _0369_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4016 _0833_/a_79_21# _0399_ _0833_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X4017 VPWR _0833_/a_79_21# _0086_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X4018 VGND _0833_/a_79_21# _0086_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4019 _0833_/a_215_47# net235 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4020 _0764_/a_81_21# _0346_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X4021 _0764_/a_299_297# _0346_ _0764_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X4022 VPWR _0764_/a_81_21# _0385_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X4023 VPWR _0373_ _0764_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4024 VGND _0764_/a_81_21# _0385_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4025 VGND _0384_ _0764_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X4026 _0764_/a_299_297# _0384_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4027 _0764_/a_384_47# _0373_ _0764_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4028 VPWR _0695_/a_80_21# _0327_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X4029 _0695_/a_80_21# _0326_ _0695_/a_472_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.31 ps=2.62 w=1 l=0.15
X4030 VPWR _0312_ _0695_/a_217_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.545 ps=5.09 w=1 l=0.15
X4031 VGND _0323_ _0695_/a_80_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.35425 ps=3.69 w=0.65 l=0.15
X4032 VGND _0695_/a_80_21# _0327_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.17225 ps=1.83 w=0.65 l=0.15
X4033 _0695_/a_300_47# _0312_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X4034 _0695_/a_217_297# _0250_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4035 _0695_/a_80_21# _0250_ _0695_/a_300_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4036 _0695_/a_472_297# _0323_ _0695_/a_217_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4037 _0695_/a_80_21# _0326_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4038 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4039 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4040 net103 clknet_1_1__leaf__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X4041 VGND clknet_1_1__leaf__0461_ net103 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X4042 net103 clknet_1_1__leaf__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4043 VPWR clknet_1_1__leaf__0461_ net103 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4044 comp0.B\[0\] _1032_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4045 _1032_/a_891_413# _1032_/a_193_47# _1032_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X4046 _1032_/a_561_413# _1032_/a_27_47# _1032_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X4047 VPWR net118 _1032_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X4048 comp0.B\[0\] _1032_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4049 _1032_/a_381_47# net202 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X4050 VGND _1032_/a_634_159# _1032_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X4051 VPWR _1032_/a_891_413# _1032_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4052 _1032_/a_466_413# _1032_/a_193_47# _1032_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4053 VPWR _1032_/a_634_159# _1032_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4054 _1032_/a_634_159# _1032_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X4055 _1032_/a_634_159# _1032_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X4056 _1032_/a_975_413# _1032_/a_193_47# _1032_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X4057 VGND _1032_/a_1059_315# _1032_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X4058 _1032_/a_193_47# _1032_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X4059 _1032_/a_891_413# _1032_/a_27_47# _1032_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4060 _1032_/a_592_47# _1032_/a_193_47# _1032_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X4061 VPWR _1032_/a_1059_315# _1032_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4062 _1032_/a_1017_47# _1032_/a_27_47# _1032_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X4063 _1032_/a_193_47# _1032_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X4064 _1032_/a_466_413# _1032_/a_27_47# _1032_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X4065 VGND _1032_/a_891_413# _1032_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4066 _1032_/a_381_47# net202 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4067 VGND net118 _1032_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4068 VGND _0218_ _0816_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4069 _0816_/a_68_297# net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4070 _0426_ _0816_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4071 VPWR _0218_ _0816_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X4072 _0426_ _0816_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X4073 _0816_/a_150_297# net67 _0816_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4074 VGND _0369_ _0747_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X4075 _0747_/a_510_47# _0371_ _0747_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X4076 _0747_/a_79_21# _0352_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X4077 VPWR _0371_ _0747_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4078 _0747_/a_79_21# net216 _0747_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X4079 _0747_/a_297_297# _0369_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4080 _0747_/a_79_21# _0352_ _0747_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X4081 VPWR _0747_/a_79_21# _0104_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X4082 VGND _0747_/a_79_21# _0104_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4083 _0747_/a_215_47# net216 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4084 VGND _0308_ _0678_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4085 _0678_/a_68_297# _0309_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4086 _0310_ _0678_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4087 VPWR _0308_ _0678_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X4088 _0310_ _0678_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X4089 _0678_/a_150_297# _0309_ _0678_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4090 VGND acc0.A\[23\] _0601_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4091 _0601_/a_68_297# net51 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4092 _0233_ _0601_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4093 VPWR acc0.A\[23\] _0601_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X4094 _0233_ _0601_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X4095 _0601_/a_150_297# net51 _0601_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4096 _0532_/a_81_21# _0198_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X4097 _0532_/a_299_297# _0198_ _0532_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X4098 VPWR _0532_/a_81_21# _0146_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X4099 VPWR net218 _0532_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4100 VGND _0532_/a_81_21# _0146_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4101 VGND _0195_ _0532_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X4102 _0532_/a_299_297# _0195_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4103 _0532_/a_384_47# net218 _0532_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4104 comp0.B\[15\] _1015_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4105 _1015_/a_891_413# _1015_/a_193_47# _1015_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X4106 _1015_/a_561_413# _1015_/a_27_47# _1015_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X4107 VPWR net101 _1015_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X4108 comp0.B\[15\] _1015_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4109 _1015_/a_381_47# _0113_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X4110 VGND _1015_/a_634_159# _1015_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X4111 VPWR _1015_/a_891_413# _1015_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4112 _1015_/a_466_413# _1015_/a_193_47# _1015_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4113 VPWR _1015_/a_634_159# _1015_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4114 _1015_/a_634_159# _1015_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X4115 _1015_/a_634_159# _1015_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X4116 _1015_/a_975_413# _1015_/a_193_47# _1015_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X4117 VGND _1015_/a_1059_315# _1015_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X4118 _1015_/a_193_47# _1015_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X4119 _1015_/a_891_413# _1015_/a_27_47# _1015_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4120 _1015_/a_592_47# _1015_/a_193_47# _1015_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X4121 VPWR _1015_/a_1059_315# _1015_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4122 _1015_/a_1017_47# _1015_/a_27_47# _1015_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X4123 _1015_/a_193_47# _1015_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X4124 _1015_/a_466_413# _1015_/a_27_47# _1015_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X4125 VGND _1015_/a_891_413# _1015_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4126 _1015_/a_381_47# _0113_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4127 VGND net101 _1015_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4128 net84 clknet_1_0__leaf__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X4129 VGND clknet_1_0__leaf__0459_ net84 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X4130 net84 clknet_1_0__leaf__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4131 VPWR clknet_1_0__leaf__0459_ net84 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4132 VPWR clknet_0__0461_ clkbuf_1_1__f__0461_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X4133 VPWR clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X4134 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4135 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4136 VPWR clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4137 VPWR clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4138 clkbuf_1_1__f__0461_/a_110_47# clknet_0__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4139 clkbuf_1_1__f__0461_/a_110_47# clknet_0__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X4140 VGND clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X4141 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4142 VGND clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4143 clkbuf_1_1__f__0461_/a_110_47# clknet_0__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4144 VGND clknet_0__0461_ clkbuf_1_1__f__0461_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4145 VGND clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4146 VPWR clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4147 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4148 VGND clknet_0__0461_ clkbuf_1_1__f__0461_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4149 VGND clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4150 VPWR clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4151 VGND clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4152 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4153 clkbuf_1_1__f__0461_/a_110_47# clknet_0__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4154 VPWR clknet_0__0461_ clkbuf_1_1__f__0461_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4155 VPWR clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4156 VPWR clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4157 VGND clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4158 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4159 VGND clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4160 VGND clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4161 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4162 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4163 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4164 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4165 VPWR clkbuf_1_1__f__0461_/a_110_47# clknet_1_1__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4166 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4167 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4168 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4169 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4170 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4171 clknet_1_1__leaf__0461_ clkbuf_1_1__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4172 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X4173 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X4174 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4175 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4176 _0515_/a_81_21# _0189_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X4177 _0515_/a_299_297# _0189_ _0515_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X4178 VPWR _0515_/a_81_21# _0154_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X4179 VPWR net181 _0515_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4180 VGND _0515_/a_81_21# _0154_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4181 VGND _0179_ _0515_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X4182 _0515_/a_299_297# _0179_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4183 _0515_/a_384_47# net181 _0515_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4184 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X4185 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X4186 net40 _0995_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4187 _0995_/a_891_413# _0995_/a_193_47# _0995_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X4188 _0995_/a_561_413# _0995_/a_27_47# _0995_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X4189 VPWR net81 _0995_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X4190 net40 _0995_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4191 _0995_/a_381_47# _0093_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X4192 VGND _0995_/a_634_159# _0995_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X4193 VPWR _0995_/a_891_413# _0995_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4194 _0995_/a_466_413# _0995_/a_193_47# _0995_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4195 VPWR _0995_/a_634_159# _0995_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4196 _0995_/a_634_159# _0995_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X4197 _0995_/a_634_159# _0995_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X4198 _0995_/a_975_413# _0995_/a_193_47# _0995_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X4199 VGND _0995_/a_1059_315# _0995_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X4200 _0995_/a_193_47# _0995_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X4201 _0995_/a_891_413# _0995_/a_27_47# _0995_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4202 _0995_/a_592_47# _0995_/a_193_47# _0995_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X4203 VPWR _0995_/a_1059_315# _0995_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4204 _0995_/a_1017_47# _0995_/a_27_47# _0995_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X4205 _0995_/a_193_47# _0995_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X4206 _0995_/a_466_413# _0995_/a_27_47# _0995_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X4207 VGND _0995_/a_891_413# _0995_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4208 _0995_/a_381_47# _0093_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4209 VGND net81 _0995_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4210 VPWR _0463_ clkbuf_0__0463_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X4211 VPWR clkbuf_0__0463_/a_110_47# clknet_0__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X4212 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4213 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4214 VPWR clkbuf_0__0463_/a_110_47# clknet_0__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4215 VPWR clkbuf_0__0463_/a_110_47# clknet_0__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4216 clkbuf_0__0463_/a_110_47# _0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4217 clkbuf_0__0463_/a_110_47# _0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X4218 VGND clkbuf_0__0463_/a_110_47# clknet_0__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X4219 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4220 VGND clkbuf_0__0463_/a_110_47# clknet_0__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4221 clkbuf_0__0463_/a_110_47# _0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4222 VGND _0463_ clkbuf_0__0463_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4223 VGND clkbuf_0__0463_/a_110_47# clknet_0__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4224 VPWR clkbuf_0__0463_/a_110_47# clknet_0__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4225 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4226 VGND _0463_ clkbuf_0__0463_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4227 VGND clkbuf_0__0463_/a_110_47# clknet_0__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4228 VPWR clkbuf_0__0463_/a_110_47# clknet_0__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4229 VGND clkbuf_0__0463_/a_110_47# clknet_0__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4230 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4231 clkbuf_0__0463_/a_110_47# _0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4232 VPWR _0463_ clkbuf_0__0463_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4233 VPWR clkbuf_0__0463_/a_110_47# clknet_0__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4234 VPWR clkbuf_0__0463_/a_110_47# clknet_0__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4235 VGND clkbuf_0__0463_/a_110_47# clknet_0__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4236 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4237 VGND clkbuf_0__0463_/a_110_47# clknet_0__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4238 VGND clkbuf_0__0463_/a_110_47# clknet_0__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4239 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4240 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4241 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4242 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4243 VPWR clkbuf_0__0463_/a_110_47# clknet_0__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4244 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4245 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4246 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4247 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4248 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4249 clknet_0__0463_ clkbuf_0__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4250 _0397_ _0780_/a_35_297# _0780_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.53 ps=5.06 w=1 l=0.15
X4251 _0397_ _0308_ _0780_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.5005 pd=2.84 as=0.1755 ps=1.84 w=0.65 l=0.15
X4252 _0780_/a_35_297# _0308_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X4253 _0780_/a_117_297# _0308_ _0780_/a_35_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.26 ps=2.52 w=1 l=0.15
X4254 VPWR _0308_ _0780_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4255 VGND _0387_ _0780_/a_35_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4256 VGND _0780_/a_35_297# _0397_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4257 _0780_/a_285_297# _0387_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4258 VPWR _0387_ _0780_/a_117_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4259 _0780_/a_285_47# _0387_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4260 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X4261 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X4262 VPWR input5/a_75_212# net5 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X4263 input5/a_75_212# A[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X4264 input5/a_75_212# A[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X4265 VGND input5/a_75_212# net5 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X4266 VPWR _0466_ _0978_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X4267 _0978_/a_27_297# _0481_ _0978_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X4268 VGND _0466_ _0978_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X4269 _0168_ _0978_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4270 _0978_/a_27_297# _0481_ _0978_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X4271 _0978_/a_109_297# net226 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4272 _0978_/a_373_47# net226 _0978_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4273 _0168_ _0978_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4274 _0978_/a_109_297# _0488_ _0978_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4275 _0978_/a_109_47# _0488_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4276 VPWR _0248_ _0384_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.53 ps=5.06 w=1 l=0.15
X4277 _0384_ _0236_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4278 _0763_/a_193_47# _0248_ _0763_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.1755 ps=1.84 w=0.65 l=0.15
X4279 _0384_ _0236_ _0763_/a_193_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4280 _0384_ _0372_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4281 _0763_/a_109_47# _0372_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4282 VPWR _0350_ _0439_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4283 _0439_ _0350_ _0832_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X4284 _0832_/a_113_47# _0438_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4285 _0439_ _0438_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4286 VPWR _0324_ _0326_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4287 _0326_ _0324_ _0694_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X4288 _0694_/a_113_47# _0325_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4289 _0326_ _0325_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4290 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X4291 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X4292 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4293 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4294 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4295 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4296 acc0.A\[31\] _1031_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4297 _1031_/a_891_413# _1031_/a_193_47# _1031_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X4298 _1031_/a_561_413# _1031_/a_27_47# _1031_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X4299 VPWR net117 _1031_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X4300 acc0.A\[31\] _1031_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4301 _1031_/a_381_47# net163 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X4302 VGND _1031_/a_634_159# _1031_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X4303 VPWR _1031_/a_891_413# _1031_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4304 _1031_/a_466_413# _1031_/a_193_47# _1031_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4305 VPWR _1031_/a_634_159# _1031_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4306 _1031_/a_634_159# _1031_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X4307 _1031_/a_634_159# _1031_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X4308 _1031_/a_975_413# _1031_/a_193_47# _1031_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X4309 VGND _1031_/a_1059_315# _1031_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X4310 _1031_/a_193_47# _1031_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X4311 _1031_/a_891_413# _1031_/a_27_47# _1031_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4312 _1031_/a_592_47# _1031_/a_193_47# _1031_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X4313 VPWR _1031_/a_1059_315# _1031_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4314 _1031_/a_1017_47# _1031_/a_27_47# _1031_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X4315 _1031_/a_193_47# _1031_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X4316 _1031_/a_466_413# _1031_/a_27_47# _1031_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X4317 VGND _1031_/a_891_413# _1031_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4318 _1031_/a_381_47# net163 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4319 VGND net117 _1031_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4320 VPWR input30/a_75_212# net30 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X4321 input30/a_75_212# B[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X4322 input30/a_75_212# B[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X4323 VGND input30/a_75_212# net30 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X4324 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4325 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4326 _0746_/a_81_21# _0346_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X4327 _0746_/a_299_297# _0346_ _0746_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X4328 VPWR _0746_/a_81_21# _0371_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X4329 VPWR _0359_ _0746_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4330 VGND _0746_/a_81_21# _0371_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4331 VGND _0370_ _0746_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X4332 _0746_/a_299_297# _0370_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4333 _0746_/a_384_47# _0359_ _0746_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4334 _0815_/a_199_47# _0290_ _0425_ VGND sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.182 ps=1.86 w=0.65 l=0.15
X4335 _0815_/a_113_297# _0401_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.545 pd=5.09 as=0 ps=0 w=1 l=0.15
X4336 _0425_ _0423_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4337 VPWR _0290_ _0815_/a_113_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4338 _0815_/a_113_297# _0423_ _0425_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X4339 VGND _0401_ _0815_/a_199_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4340 _0677_/a_377_297# acc0.A\[17\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=2.42 as=0 ps=0 w=1 l=0.15
X4341 _0677_/a_47_47# net44 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X4342 _0677_/a_129_47# net44 _0677_/a_47_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.72 as=0.169 ps=1.82 w=0.65 l=0.15
X4343 _0677_/a_285_47# net44 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X4344 _0309_ _0677_/a_47_47# _0677_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X4345 VGND acc0.A\[17\] _0677_/a_129_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4346 VPWR acc0.A\[17\] _0677_/a_47_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4347 VPWR _0677_/a_47_47# _0309_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.33 ps=2.66 w=1 l=0.15
X4348 _0309_ net44 _0677_/a_377_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4349 _0677_/a_285_47# acc0.A\[17\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4350 _0600_/a_103_199# _0231_ _0600_/a_253_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.39 ps=3.8 w=0.65 l=0.15
X4351 VPWR _0600_/a_103_199# _0232_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.36 ps=2.72 w=1 l=0.15
X4352 _0600_/a_337_297# _0223_ _0600_/a_253_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.27 ps=2.54 w=1 l=0.15
X4353 _0600_/a_103_199# _0230_ _0600_/a_337_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.425 pd=2.85 as=0 ps=0 w=1 l=0.15
X4354 _0600_/a_253_297# _0225_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4355 VPWR _0231_ _0600_/a_103_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4356 VGND _0600_/a_103_199# _0232_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.234 ps=2.02 w=0.65 l=0.15
X4357 _0600_/a_253_47# _0225_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4358 _0600_/a_253_47# _0230_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4359 VGND _0223_ _0600_/a_253_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4360 VPWR net9 _0531_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X4361 _0531_/a_27_297# _0182_ _0531_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X4362 VGND net9 _0531_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X4363 _0198_ _0531_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4364 _0531_/a_27_297# _0182_ _0531_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X4365 _0531_/a_109_297# _0180_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4366 _0531_/a_373_47# _0180_ _0531_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4367 _0198_ _0531_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4368 _0531_/a_109_297# net175 _0531_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4369 _0531_/a_109_47# net175 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4370 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4371 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4372 acc0.A\[0\] _1014_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4373 _1014_/a_891_413# _1014_/a_193_47# _1014_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X4374 _1014_/a_561_413# _1014_/a_27_47# _1014_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X4375 VPWR net100 _1014_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X4376 acc0.A\[0\] _1014_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4377 _1014_/a_381_47# _0112_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X4378 VGND _1014_/a_634_159# _1014_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X4379 VPWR _1014_/a_891_413# _1014_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4380 _1014_/a_466_413# _1014_/a_193_47# _1014_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4381 VPWR _1014_/a_634_159# _1014_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4382 _1014_/a_634_159# _1014_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X4383 _1014_/a_634_159# _1014_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X4384 _1014_/a_975_413# _1014_/a_193_47# _1014_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X4385 VGND _1014_/a_1059_315# _1014_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X4386 _1014_/a_193_47# _1014_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X4387 _1014_/a_891_413# _1014_/a_27_47# _1014_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4388 _1014_/a_592_47# _1014_/a_193_47# _1014_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X4389 VPWR _1014_/a_1059_315# _1014_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4390 _1014_/a_1017_47# _1014_/a_27_47# _1014_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X4391 _1014_/a_193_47# _1014_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X4392 _1014_/a_466_413# _1014_/a_27_47# _1014_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X4393 VGND _1014_/a_891_413# _1014_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4394 _1014_/a_381_47# _0112_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4395 VGND net100 _1014_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4396 VGND _0350_ _0729_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4397 _0729_/a_68_297# net242 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4398 _0358_ _0729_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4399 VPWR _0350_ _0729_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X4400 _0358_ _0729_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X4401 _0729_/a_150_297# net242 _0729_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4402 net141 clknet_1_1__leaf__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X4403 VGND clknet_1_1__leaf__0465_ net141 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X4404 net141 clknet_1_1__leaf__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4405 VPWR clknet_1_1__leaf__0465_ net141 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4406 VPWR clknet_0__0460_ clkbuf_1_1__f__0460_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X4407 VPWR clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X4408 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4409 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4410 VPWR clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4411 VPWR clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4412 clkbuf_1_1__f__0460_/a_110_47# clknet_0__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4413 clkbuf_1_1__f__0460_/a_110_47# clknet_0__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X4414 VGND clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X4415 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4416 VGND clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4417 clkbuf_1_1__f__0460_/a_110_47# clknet_0__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4418 VGND clknet_0__0460_ clkbuf_1_1__f__0460_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4419 VGND clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4420 VPWR clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4421 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4422 VGND clknet_0__0460_ clkbuf_1_1__f__0460_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4423 VGND clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4424 VPWR clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4425 VGND clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4426 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4427 clkbuf_1_1__f__0460_/a_110_47# clknet_0__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4428 VPWR clknet_0__0460_ clkbuf_1_1__f__0460_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4429 VPWR clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4430 VPWR clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4431 VGND clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4432 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4433 VGND clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4434 VGND clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4435 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4436 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4437 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4438 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4439 VPWR clkbuf_1_1__f__0460_/a_110_47# clknet_1_1__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4440 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4441 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4442 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4443 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4444 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4445 clknet_1_1__leaf__0460_ clkbuf_1_1__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4446 net71 clknet_1_0__leaf__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X4447 VGND clknet_1_0__leaf__0458_ net71 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X4448 net71 clknet_1_0__leaf__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4449 VPWR clknet_1_0__leaf__0458_ net71 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4450 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4451 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4452 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X4453 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X4454 net88 clknet_1_0__leaf__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X4455 VGND clknet_1_0__leaf__0460_ net88 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X4456 net88 clknet_1_0__leaf__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4457 VPWR clknet_1_0__leaf__0460_ net88 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4458 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4459 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4460 VPWR net2 _0514_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X4461 _0514_/a_27_297# _0186_ _0514_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X4462 VGND net2 _0514_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X4463 _0189_ _0514_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4464 _0514_/a_27_297# _0186_ _0514_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X4465 _0514_/a_109_297# _0181_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4466 _0514_/a_373_47# _0181_ _0514_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4467 _0189_ _0514_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4468 _0514_/a_109_297# acc0.A\[10\] _0514_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4469 _0514_/a_109_47# acc0.A\[10\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4470 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4471 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4472 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4473 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4474 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4475 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4476 net122 clknet_1_1__leaf__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X4477 VGND clknet_1_1__leaf__0463_ net122 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X4478 net122 clknet_1_1__leaf__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4479 VPWR clknet_1_1__leaf__0463_ net122 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4480 net136 clknet_1_0__leaf__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X4481 VGND clknet_1_0__leaf__0464_ net136 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X4482 net136 clknet_1_0__leaf__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4483 VPWR clknet_1_0__leaf__0464_ net136 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4484 net39 _0994_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4485 _0994_/a_891_413# _0994_/a_193_47# _0994_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X4486 _0994_/a_561_413# _0994_/a_27_47# _0994_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X4487 VPWR net80 _0994_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X4488 net39 _0994_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4489 _0994_/a_381_47# _0092_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X4490 VGND _0994_/a_634_159# _0994_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X4491 VPWR _0994_/a_891_413# _0994_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4492 _0994_/a_466_413# _0994_/a_193_47# _0994_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4493 VPWR _0994_/a_634_159# _0994_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4494 _0994_/a_634_159# _0994_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X4495 _0994_/a_634_159# _0994_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X4496 _0994_/a_975_413# _0994_/a_193_47# _0994_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X4497 VGND _0994_/a_1059_315# _0994_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X4498 _0994_/a_193_47# _0994_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X4499 _0994_/a_891_413# _0994_/a_27_47# _0994_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4500 _0994_/a_592_47# _0994_/a_193_47# _0994_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X4501 VPWR _0994_/a_1059_315# _0994_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4502 _0994_/a_1017_47# _0994_/a_27_47# _0994_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X4503 _0994_/a_193_47# _0994_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X4504 _0994_/a_466_413# _0994_/a_27_47# _0994_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X4505 VGND _0994_/a_891_413# _0994_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4506 _0994_/a_381_47# _0092_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4507 VGND net80 _0994_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4508 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4509 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4510 VPWR _0462_ clkbuf_0__0462_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X4511 VPWR clkbuf_0__0462_/a_110_47# clknet_0__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X4512 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4513 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4514 VPWR clkbuf_0__0462_/a_110_47# clknet_0__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4515 VPWR clkbuf_0__0462_/a_110_47# clknet_0__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4516 clkbuf_0__0462_/a_110_47# _0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4517 clkbuf_0__0462_/a_110_47# _0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X4518 VGND clkbuf_0__0462_/a_110_47# clknet_0__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X4519 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4520 VGND clkbuf_0__0462_/a_110_47# clknet_0__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4521 clkbuf_0__0462_/a_110_47# _0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4522 VGND _0462_ clkbuf_0__0462_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4523 VGND clkbuf_0__0462_/a_110_47# clknet_0__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4524 VPWR clkbuf_0__0462_/a_110_47# clknet_0__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4525 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4526 VGND _0462_ clkbuf_0__0462_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4527 VGND clkbuf_0__0462_/a_110_47# clknet_0__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4528 VPWR clkbuf_0__0462_/a_110_47# clknet_0__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4529 VGND clkbuf_0__0462_/a_110_47# clknet_0__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4530 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4531 clkbuf_0__0462_/a_110_47# _0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4532 VPWR _0462_ clkbuf_0__0462_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4533 VPWR clkbuf_0__0462_/a_110_47# clknet_0__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4534 VPWR clkbuf_0__0462_/a_110_47# clknet_0__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4535 VGND clkbuf_0__0462_/a_110_47# clknet_0__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4536 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4537 VGND clkbuf_0__0462_/a_110_47# clknet_0__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4538 VGND clkbuf_0__0462_/a_110_47# clknet_0__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4539 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4540 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4541 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4542 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4543 VPWR clkbuf_0__0462_/a_110_47# clknet_0__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4544 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4545 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4546 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4547 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4548 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4549 clknet_0__0462_ clkbuf_0__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4550 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X4551 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X4552 VPWR input6/a_75_212# net6 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X4553 input6/a_75_212# A[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X4554 input6/a_75_212# A[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X4555 VGND input6/a_75_212# net6 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X4556 VPWR _0977_/a_75_212# _0167_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X4557 _0977_/a_75_212# _0489_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X4558 _0977_/a_75_212# _0489_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X4559 VGND _0977_/a_75_212# _0167_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X4560 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4561 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4562 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4563 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4564 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4565 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4566 _0438_ _0831_/a_35_297# _0831_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.53 ps=5.06 w=1 l=0.15
X4567 _0438_ _0434_ _0831_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.5005 pd=2.84 as=0.1755 ps=1.84 w=0.65 l=0.15
X4568 _0831_/a_35_297# _0434_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X4569 _0831_/a_117_297# _0434_ _0831_/a_35_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.26 ps=2.52 w=1 l=0.15
X4570 VPWR _0434_ _0831_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4571 VGND _0253_ _0831_/a_35_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4572 VGND _0831_/a_35_297# _0438_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4573 _0831_/a_285_297# _0253_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4574 VPWR _0253_ _0831_/a_117_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4575 _0831_/a_285_47# _0253_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4576 VGND _0369_ _0762_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X4577 _0762_/a_510_47# _0383_ _0762_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X4578 _0762_/a_79_21# _0352_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X4579 VPWR _0383_ _0762_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4580 _0762_/a_79_21# net213 _0762_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X4581 _0762_/a_297_297# _0369_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4582 _0762_/a_79_21# _0352_ _0762_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X4583 VPWR _0762_/a_79_21# _0101_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X4584 VGND _0762_/a_79_21# _0101_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4585 _0762_/a_215_47# net213 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4586 VGND acc0.A\[24\] _0693_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4587 _0693_/a_68_297# net52 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4588 _0325_ _0693_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4589 VPWR acc0.A\[24\] _0693_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X4590 _0325_ _0693_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X4591 _0693_/a_150_297# net52 _0693_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4592 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4593 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4594 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X4595 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X4596 acc0.A\[30\] _1030_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4597 _1030_/a_891_413# _1030_/a_193_47# _1030_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X4598 _1030_/a_561_413# _1030_/a_27_47# _1030_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X4599 VPWR net116 _1030_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X4600 acc0.A\[30\] _1030_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4601 _1030_/a_381_47# net209 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X4602 VGND _1030_/a_634_159# _1030_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X4603 VPWR _1030_/a_891_413# _1030_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4604 _1030_/a_466_413# _1030_/a_193_47# _1030_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4605 VPWR _1030_/a_634_159# _1030_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4606 _1030_/a_634_159# _1030_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X4607 _1030_/a_634_159# _1030_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X4608 _1030_/a_975_413# _1030_/a_193_47# _1030_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X4609 VGND _1030_/a_1059_315# _1030_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X4610 _1030_/a_193_47# _1030_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X4611 _1030_/a_891_413# _1030_/a_27_47# _1030_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4612 _1030_/a_592_47# _1030_/a_193_47# _1030_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X4613 VPWR _1030_/a_1059_315# _1030_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4614 _1030_/a_1017_47# _1030_/a_27_47# _1030_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X4615 _1030_/a_193_47# _1030_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X4616 _1030_/a_466_413# _1030_/a_27_47# _1030_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X4617 VGND _1030_/a_891_413# _1030_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4618 _1030_/a_381_47# net209 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4619 VGND net116 _1030_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4620 VPWR input20/a_75_212# net20 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X4621 input20/a_75_212# B[12] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X4622 input20/a_75_212# B[12] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X4623 VGND input20/a_75_212# net20 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X4624 VPWR input31/a_75_212# net31 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X4625 input31/a_75_212# B[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X4626 input31/a_75_212# B[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X4627 VGND input31/a_75_212# net31 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X4628 VPWR _0423_ _0814_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2415 ps=2.83 w=0.42 l=0.15
X4629 VPWR _0401_ _0814_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4630 _0814_/a_181_47# _0290_ _0814_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0882 pd=1.26 as=0.0882 ps=1.26 w=0.42 l=0.15
X4631 VGND _0401_ _0814_/a_181_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4632 _0814_/a_27_47# _0290_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4633 _0424_ _0814_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4634 _0424_ _0814_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4635 _0814_/a_109_47# _0423_ _0814_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4636 VPWR _0250_ _0370_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.53 ps=5.06 w=1 l=0.15
X4637 _0370_ _0326_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4638 _0745_/a_193_47# _0250_ _0745_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.1755 ps=1.84 w=0.65 l=0.15
X4639 _0370_ _0326_ _0745_/a_193_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4640 _0370_ _0312_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4641 _0745_/a_109_47# _0312_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4642 VPWR _0306_ _0308_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4643 _0308_ _0306_ _0676_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X4644 _0676_/a_113_47# _0307_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4645 _0308_ _0307_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4646 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4647 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4648 _0530_/a_81_21# _0197_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X4649 _0530_/a_299_297# _0197_ _0530_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X4650 VPWR _0530_/a_81_21# _0147_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X4651 VPWR net175 _0530_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4652 VGND _0530_/a_81_21# _0147_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4653 VGND _0195_ _0530_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X4654 _0530_/a_299_297# _0195_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4655 _0530_/a_384_47# net175 _0530_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4656 net60 _1013_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4657 _1013_/a_891_413# _1013_/a_193_47# _1013_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X4658 _1013_/a_561_413# _1013_/a_27_47# _1013_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X4659 VPWR net99 _1013_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X4660 net60 _1013_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4661 _1013_/a_381_47# _0111_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X4662 VGND _1013_/a_634_159# _1013_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X4663 VPWR _1013_/a_891_413# _1013_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4664 _1013_/a_466_413# _1013_/a_193_47# _1013_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4665 VPWR _1013_/a_634_159# _1013_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4666 _1013_/a_634_159# _1013_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X4667 _1013_/a_634_159# _1013_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X4668 _1013_/a_975_413# _1013_/a_193_47# _1013_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X4669 VGND _1013_/a_1059_315# _1013_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X4670 _1013_/a_193_47# _1013_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X4671 _1013_/a_891_413# _1013_/a_27_47# _1013_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4672 _1013_/a_592_47# _1013_/a_193_47# _1013_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X4673 VPWR _1013_/a_1059_315# _1013_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4674 _1013_/a_1017_47# _1013_/a_27_47# _1013_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X4675 _1013_/a_193_47# _1013_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X4676 _1013_/a_466_413# _1013_/a_27_47# _1013_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X4677 VGND _1013_/a_891_413# _1013_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4678 _1013_/a_381_47# _0111_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4679 VGND net99 _1013_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4680 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4681 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4682 VPWR _0356_ _0728_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4683 _0357_ _0728_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X4684 VGND _0356_ _0728_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4685 _0728_/a_59_75# _0333_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4686 _0357_ _0728_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X4687 _0728_/a_145_75# _0333_ _0728_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X4688 VGND acc0.A\[8\] _0659_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4689 _0659_/a_68_297# net66 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4690 _0291_ _0659_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4691 VPWR acc0.A\[8\] _0659_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X4692 _0291_ _0659_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X4693 _0659_/a_150_297# net66 _0659_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4694 _0513_/a_81_21# _0188_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X4695 _0513_/a_299_297# _0188_ _0513_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X4696 VPWR _0513_/a_81_21# _0155_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X4697 VPWR net188 _0513_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4698 VGND _0513_/a_81_21# _0155_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4699 VGND _0179_ _0513_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X4700 _0513_/a_299_297# _0179_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4701 _0513_/a_384_47# net188 _0513_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4702 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4703 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4704 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4705 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4706 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4707 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4708 net38 _0993_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4709 _0993_/a_891_413# _0993_/a_193_47# _0993_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X4710 _0993_/a_561_413# _0993_/a_27_47# _0993_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X4711 VPWR net79 _0993_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X4712 net38 _0993_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4713 _0993_/a_381_47# _0091_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X4714 VGND _0993_/a_634_159# _0993_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X4715 VPWR _0993_/a_891_413# _0993_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4716 _0993_/a_466_413# _0993_/a_193_47# _0993_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4717 VPWR _0993_/a_634_159# _0993_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4718 _0993_/a_634_159# _0993_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X4719 _0993_/a_634_159# _0993_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X4720 _0993_/a_975_413# _0993_/a_193_47# _0993_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X4721 VGND _0993_/a_1059_315# _0993_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X4722 _0993_/a_193_47# _0993_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X4723 _0993_/a_891_413# _0993_/a_27_47# _0993_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4724 _0993_/a_592_47# _0993_/a_193_47# _0993_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X4725 VPWR _0993_/a_1059_315# _0993_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4726 _0993_/a_1017_47# _0993_/a_27_47# _0993_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X4727 _0993_/a_193_47# _0993_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X4728 _0993_/a_466_413# _0993_/a_27_47# _0993_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X4729 VGND _0993_/a_891_413# _0993_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4730 _0993_/a_381_47# _0091_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4731 VGND net79 _0993_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4732 VPWR _0461_ clkbuf_0__0461_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X4733 VPWR clkbuf_0__0461_/a_110_47# clknet_0__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X4734 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4735 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4736 VPWR clkbuf_0__0461_/a_110_47# clknet_0__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4737 VPWR clkbuf_0__0461_/a_110_47# clknet_0__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4738 clkbuf_0__0461_/a_110_47# _0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4739 clkbuf_0__0461_/a_110_47# _0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X4740 VGND clkbuf_0__0461_/a_110_47# clknet_0__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X4741 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4742 VGND clkbuf_0__0461_/a_110_47# clknet_0__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4743 clkbuf_0__0461_/a_110_47# _0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4744 VGND _0461_ clkbuf_0__0461_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4745 VGND clkbuf_0__0461_/a_110_47# clknet_0__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4746 VPWR clkbuf_0__0461_/a_110_47# clknet_0__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4747 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4748 VGND _0461_ clkbuf_0__0461_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4749 VGND clkbuf_0__0461_/a_110_47# clknet_0__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4750 VPWR clkbuf_0__0461_/a_110_47# clknet_0__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4751 VGND clkbuf_0__0461_/a_110_47# clknet_0__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4752 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4753 clkbuf_0__0461_/a_110_47# _0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4754 VPWR _0461_ clkbuf_0__0461_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4755 VPWR clkbuf_0__0461_/a_110_47# clknet_0__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4756 VPWR clkbuf_0__0461_/a_110_47# clknet_0__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4757 VGND clkbuf_0__0461_/a_110_47# clknet_0__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4758 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4759 VGND clkbuf_0__0461_/a_110_47# clknet_0__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4760 VGND clkbuf_0__0461_/a_110_47# clknet_0__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4761 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4762 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4763 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4764 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4765 VPWR clkbuf_0__0461_/a_110_47# clknet_0__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4766 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4767 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4768 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4769 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4770 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4771 clknet_0__0461_ clkbuf_0__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4772 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4773 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4774 VPWR input7/a_75_212# net7 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X4775 input7/a_75_212# A[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X4776 input7/a_75_212# A[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X4777 VGND input7/a_75_212# net7 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X4778 VPWR _0976_/a_505_21# _0976_/a_535_374# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4779 _0976_/a_505_21# control0.count\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X4780 _0976_/a_218_374# control0.count\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X4781 VGND _0976_/a_505_21# _0976_/a_439_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4782 _0976_/a_76_199# _0488_ _0976_/a_218_374# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X4783 _0976_/a_505_21# control0.count\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X4784 _0976_/a_439_47# _0488_ _0976_/a_76_199# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X4785 _0976_/a_535_374# _0466_ _0976_/a_76_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X4786 _0976_/a_76_199# _0466_ _0976_/a_218_47# VGND sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X4787 _0976_/a_218_47# control0.count\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X4788 VPWR _0976_/a_76_199# _0489_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X4789 VGND _0976_/a_76_199# _0489_ VGND sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
X4790 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X4791 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X4792 VGND _0369_ _0830_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X4793 _0830_/a_510_47# _0437_ _0830_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X4794 _0830_/a_79_21# _0399_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X4795 VPWR _0437_ _0830_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4796 _0830_/a_79_21# net212 _0830_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X4797 _0830_/a_297_297# _0369_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4798 _0830_/a_79_21# _0399_ _0830_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X4799 VPWR _0830_/a_79_21# _0087_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X4800 VGND _0830_/a_79_21# _0087_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4801 _0830_/a_215_47# net212 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4802 VPWR _0219_ _0383_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4803 _0383_ _0219_ _0761_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X4804 _0761_/a_113_47# _0382_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4805 _0383_ _0382_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4806 VPWR acc0.A\[24\] _0324_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4807 _0324_ acc0.A\[24\] _0692_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X4808 _0692_/a_113_47# net52 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4809 _0324_ net52 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4810 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X4811 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X4812 VPWR _0959_/a_80_21# _0160_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X4813 _0959_/a_80_21# _0477_ _0959_/a_472_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.31 ps=2.62 w=1 l=0.15
X4814 VPWR _0467_ _0959_/a_217_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.545 ps=5.09 w=1 l=0.15
X4815 VGND _0470_ _0959_/a_80_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.35425 ps=3.69 w=0.65 l=0.15
X4816 VGND _0959_/a_80_21# _0160_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.17225 ps=1.83 w=0.65 l=0.15
X4817 _0959_/a_300_47# _0467_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X4818 _0959_/a_217_297# net33 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4819 _0959_/a_80_21# net33 _0959_/a_300_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4820 _0959_/a_472_297# _0470_ _0959_/a_217_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4821 _0959_/a_80_21# _0477_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4822 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X4823 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X4824 net95 clknet_1_1__leaf__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X4825 VGND clknet_1_1__leaf__0460_ net95 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X4826 net95 clknet_1_1__leaf__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4827 VPWR clknet_1_1__leaf__0460_ net95 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4828 VPWR input10/a_75_212# net10 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X4829 input10/a_75_212# A[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X4830 input10/a_75_212# A[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X4831 VGND input10/a_75_212# net10 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X4832 VPWR input21/a_75_212# net21 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X4833 input21/a_75_212# B[13] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X4834 input21/a_75_212# B[13] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X4835 VGND input21/a_75_212# net21 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X4836 VPWR input32/a_75_212# net32 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X4837 input32/a_75_212# B[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X4838 input32/a_75_212# B[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X4839 VGND input32/a_75_212# net32 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X4840 VPWR _0288_ _0813_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X4841 VGND _0288_ _0423_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X4842 _0813_/a_109_297# _0289_ _0423_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X4843 _0423_ _0289_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4844 VPWR _0350_ _0744_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X4845 VGND _0744_/a_27_47# _0369_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X4846 VGND _0744_/a_27_47# _0369_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4847 _0369_ _0744_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X4848 _0369_ _0744_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4849 VGND _0350_ _0744_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X4850 VPWR _0744_/a_27_47# _0369_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4851 _0369_ _0744_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4852 _0369_ _0744_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4853 VPWR _0744_/a_27_47# _0369_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4854 VGND acc0.A\[16\] _0675_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4855 _0675_/a_68_297# net43 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4856 _0307_ _0675_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4857 VPWR acc0.A\[16\] _0675_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X4858 _0307_ _0675_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X4859 _0675_/a_150_297# net43 _0675_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4860 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X4861 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X4862 net59 _1012_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4863 _1012_/a_891_413# _1012_/a_193_47# _1012_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X4864 _1012_/a_561_413# _1012_/a_27_47# _1012_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X4865 VPWR net98 _1012_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X4866 net59 _1012_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4867 _1012_/a_381_47# _0110_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X4868 VGND _1012_/a_634_159# _1012_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X4869 VPWR _1012_/a_891_413# _1012_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4870 _1012_/a_466_413# _1012_/a_193_47# _1012_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4871 VPWR _1012_/a_634_159# _1012_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4872 _1012_/a_634_159# _1012_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X4873 _1012_/a_634_159# _1012_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X4874 _1012_/a_975_413# _1012_/a_193_47# _1012_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X4875 VGND _1012_/a_1059_315# _1012_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X4876 _1012_/a_193_47# _1012_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X4877 _1012_/a_891_413# _1012_/a_27_47# _1012_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4878 _1012_/a_592_47# _1012_/a_193_47# _1012_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X4879 VPWR _1012_/a_1059_315# _1012_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4880 _1012_/a_1017_47# _1012_/a_27_47# _1012_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X4881 _1012_/a_193_47# _1012_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X4882 _1012_/a_466_413# _1012_/a_27_47# _1012_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X4883 VGND _1012_/a_891_413# _1012_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4884 _1012_/a_381_47# _0110_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4885 VGND net98 _1012_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4886 _0356_ _0327_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X4887 VPWR _0332_ _0356_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.165 ps=1.33 w=1 l=0.15
X4888 VPWR _0329_ _0356_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4889 _0727_/a_193_47# _0329_ _0727_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4890 _0356_ _0332_ _0727_/a_277_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.10725 ps=0.98 w=0.65 l=0.15
X4891 _0727_/a_277_47# _0327_ _0727_/a_193_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X4892 _0356_ _0330_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X4893 _0727_/a_109_47# _0330_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X4894 VPWR acc0.A\[8\] _0290_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4895 _0290_ acc0.A\[8\] _0658_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X4896 _0658_/a_113_47# net66 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4897 _0290_ net66 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4898 VPWR acc0.A\[28\] _0221_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4899 _0221_ acc0.A\[28\] _0589_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X4900 _0589_/a_113_47# net56 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4901 _0221_ net56 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4902 VPWR net3 _0512_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X4903 _0512_/a_27_297# _0186_ _0512_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X4904 VGND net3 _0512_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X4905 _0188_ _0512_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4906 _0512_/a_27_297# _0186_ _0512_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X4907 _0512_/a_109_297# _0181_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4908 _0512_/a_373_47# _0181_ _0512_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4909 _0188_ _0512_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4910 _0512_/a_109_297# acc0.A\[11\] _0512_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4911 _0512_/a_109_47# acc0.A\[11\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4912 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4913 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4914 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4915 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X4916 net37 _0992_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X4917 _0992_/a_891_413# _0992_/a_193_47# _0992_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X4918 _0992_/a_561_413# _0992_/a_27_47# _0992_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X4919 VPWR net78 _0992_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X4920 net37 _0992_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X4921 _0992_/a_381_47# _0090_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X4922 VGND _0992_/a_634_159# _0992_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X4923 VPWR _0992_/a_891_413# _0992_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X4924 _0992_/a_466_413# _0992_/a_193_47# _0992_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4925 VPWR _0992_/a_634_159# _0992_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4926 _0992_/a_634_159# _0992_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X4927 _0992_/a_634_159# _0992_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X4928 _0992_/a_975_413# _0992_/a_193_47# _0992_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X4929 VGND _0992_/a_1059_315# _0992_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X4930 _0992_/a_193_47# _0992_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X4931 _0992_/a_891_413# _0992_/a_27_47# _0992_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4932 _0992_/a_592_47# _0992_/a_193_47# _0992_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X4933 VPWR _0992_/a_1059_315# _0992_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4934 _0992_/a_1017_47# _0992_/a_27_47# _0992_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X4935 _0992_/a_193_47# _0992_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X4936 _0992_/a_466_413# _0992_/a_27_47# _0992_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X4937 VGND _0992_/a_891_413# _0992_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X4938 _0992_/a_381_47# _0090_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4939 VGND net78 _0992_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X4940 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X4941 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X4942 VPWR _0460_ clkbuf_0__0460_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X4943 VPWR clkbuf_0__0460_/a_110_47# clknet_0__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X4944 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4945 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4946 VPWR clkbuf_0__0460_/a_110_47# clknet_0__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4947 VPWR clkbuf_0__0460_/a_110_47# clknet_0__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4948 clkbuf_0__0460_/a_110_47# _0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4949 clkbuf_0__0460_/a_110_47# _0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X4950 VGND clkbuf_0__0460_/a_110_47# clknet_0__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X4951 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4952 VGND clkbuf_0__0460_/a_110_47# clknet_0__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4953 clkbuf_0__0460_/a_110_47# _0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4954 VGND _0460_ clkbuf_0__0460_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4955 VGND clkbuf_0__0460_/a_110_47# clknet_0__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4956 VPWR clkbuf_0__0460_/a_110_47# clknet_0__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4957 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4958 VGND _0460_ clkbuf_0__0460_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4959 VGND clkbuf_0__0460_/a_110_47# clknet_0__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4960 VPWR clkbuf_0__0460_/a_110_47# clknet_0__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4961 VGND clkbuf_0__0460_/a_110_47# clknet_0__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4962 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4963 clkbuf_0__0460_/a_110_47# _0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4964 VPWR _0460_ clkbuf_0__0460_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4965 VPWR clkbuf_0__0460_/a_110_47# clknet_0__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4966 VPWR clkbuf_0__0460_/a_110_47# clknet_0__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4967 VGND clkbuf_0__0460_/a_110_47# clknet_0__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4968 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4969 VGND clkbuf_0__0460_/a_110_47# clknet_0__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4970 VGND clkbuf_0__0460_/a_110_47# clknet_0__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4971 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4972 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4973 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4974 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4975 VPWR clkbuf_0__0460_/a_110_47# clknet_0__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4976 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4977 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4978 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4979 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4980 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4981 clknet_0__0460_ clkbuf_0__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4982 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X4983 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X4984 net127 clknet_1_0__leaf__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X4985 VGND clknet_1_0__leaf__0463_ net127 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X4986 net127 clknet_1_0__leaf__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X4987 VPWR clknet_1_0__leaf__0463_ net127 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X4988 VPWR input8/a_75_212# net8 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X4989 input8/a_75_212# A[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X4990 input8/a_75_212# A[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X4991 VGND input8/a_75_212# net8 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X4992 VPWR _0486_ _0975_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4993 _0488_ _0975_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X4994 VGND _0486_ _0975_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X4995 _0975_/a_59_75# control0.state\[2\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X4996 _0488_ _0975_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X4997 _0975_/a_145_75# control0.state\[2\] _0975_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X4998 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X4999 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5000 _0760_/a_377_297# _0237_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=2.42 as=0 ps=0 w=1 l=0.15
X5001 _0760_/a_47_47# _0381_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X5002 _0760_/a_129_47# _0381_ _0760_/a_47_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.72 as=0.169 ps=1.82 w=0.65 l=0.15
X5003 _0760_/a_285_47# _0381_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X5004 _0382_ _0760_/a_47_47# _0760_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X5005 VGND _0237_ _0760_/a_129_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5006 VPWR _0237_ _0760_/a_47_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5007 VPWR _0760_/a_47_47# _0382_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.33 ps=2.66 w=1 l=0.15
X5008 _0382_ _0381_ _0760_/a_377_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5009 _0760_/a_285_47# _0237_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5010 VGND _0315_ _0691_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X5011 _0691_/a_68_297# _0322_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5012 _0323_ _0691_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5013 VPWR _0315_ _0691_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X5014 _0323_ _0691_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X5015 _0691_/a_150_297# _0322_ _0691_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5016 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5017 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5018 _0958_/a_27_47# _0476_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X5019 _0958_/a_197_47# _0471_ _0958_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X5020 _0477_ _0958_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.31245 ps=1.68 w=1 l=0.15
X5021 _0958_/a_303_47# _0476_ _0958_/a_197_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X5022 _0958_/a_27_47# control0.state\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.1092 ps=1.36 w=0.42 l=0.15
X5023 VPWR _0468_ _0958_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.31245 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X5024 VGND _0468_ _0958_/a_303_47# VGND sky130_fd_pr__nfet_01v8 ad=0.19627 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X5025 VPWR _0471_ _0958_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X5026 _0477_ _0958_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.19627 ps=1.33 w=0.65 l=0.15
X5027 _0958_/a_109_47# control0.state\[1\] _0958_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X5028 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5029 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5030 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5031 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5032 _0743_/a_240_47# net237 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X5033 _0105_ _0743_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X5034 VGND _0219_ _0743_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5035 _0743_/a_51_297# _0368_ _0743_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X5036 _0743_/a_149_47# _0345_ _0743_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X5037 _0743_/a_240_47# _0367_ _0743_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5038 VPWR _0219_ _0743_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X5039 _0105_ _0743_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X5040 _0743_/a_149_47# _0368_ _0743_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5041 _0743_/a_245_297# _0367_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5042 VPWR _0345_ _0743_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5043 _0743_/a_512_297# net237 _0743_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5044 VPWR input11/a_75_212# net11 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5045 input11/a_75_212# A[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5046 input11/a_75_212# A[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5047 VGND input11/a_75_212# net11 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5048 VPWR input22/a_75_212# net22 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5049 input22/a_75_212# B[14] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5050 input22/a_75_212# B[14] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5051 VGND input22/a_75_212# net22 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5052 VPWR input33/a_75_212# net33 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5053 input33/a_75_212# init VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5054 input33/a_75_212# init VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5055 VGND input33/a_75_212# net33 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5056 VGND _0369_ _0812_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X5057 _0812_/a_510_47# _0422_ _0812_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X5058 _0812_/a_79_21# _0399_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X5059 VPWR _0422_ _0812_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5060 _0812_/a_79_21# net217 _0812_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X5061 _0812_/a_297_297# _0369_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5062 _0812_/a_79_21# _0399_ _0812_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X5063 VPWR _0812_/a_79_21# _0090_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5064 VGND _0812_/a_79_21# _0090_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5065 _0812_/a_215_47# net217 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5066 VPWR acc0.A\[16\] _0306_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5067 _0306_ acc0.A\[16\] _0674_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X5068 _0674_/a_113_47# net43 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5069 _0306_ net43 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5070 VPWR clknet_0_clk clkbuf_1_0__f_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X5071 VPWR clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X5072 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5073 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5074 VPWR clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5075 VPWR clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5076 clkbuf_1_0__f_clk/a_110_47# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5077 clkbuf_1_0__f_clk/a_110_47# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X5078 VGND clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X5079 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5080 VGND clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5081 clkbuf_1_0__f_clk/a_110_47# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5082 VGND clknet_0_clk clkbuf_1_0__f_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5083 VGND clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5084 VPWR clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5085 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5086 VGND clknet_0_clk clkbuf_1_0__f_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5087 VGND clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5088 VPWR clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5089 VGND clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5090 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5091 clkbuf_1_0__f_clk/a_110_47# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5092 VPWR clknet_0_clk clkbuf_1_0__f_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5093 VPWR clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5094 VPWR clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5095 VGND clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5096 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5097 VGND clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5098 VGND clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5099 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5100 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5101 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5102 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5103 VPWR clkbuf_1_0__f_clk/a_110_47# clknet_1_0__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5104 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5105 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5106 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5107 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5108 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5109 clknet_1_0__leaf_clk clkbuf_1_0__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5110 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5111 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5112 net99 clknet_1_1__leaf__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X5113 VGND clknet_1_1__leaf__0461_ net99 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X5114 net99 clknet_1_1__leaf__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5115 VPWR clknet_1_1__leaf__0461_ net99 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5116 net57 _1011_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5117 _1011_/a_891_413# _1011_/a_193_47# _1011_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X5118 _1011_/a_561_413# _1011_/a_27_47# _1011_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X5119 VPWR net97 _1011_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X5120 net57 _1011_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5121 _1011_/a_381_47# _0109_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X5122 VGND _1011_/a_634_159# _1011_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X5123 VPWR _1011_/a_891_413# _1011_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5124 _1011_/a_466_413# _1011_/a_193_47# _1011_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5125 VPWR _1011_/a_634_159# _1011_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5126 _1011_/a_634_159# _1011_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X5127 _1011_/a_634_159# _1011_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X5128 _1011_/a_975_413# _1011_/a_193_47# _1011_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X5129 VGND _1011_/a_1059_315# _1011_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X5130 _1011_/a_193_47# _1011_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X5131 _1011_/a_891_413# _1011_/a_27_47# _1011_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5132 _1011_/a_592_47# _1011_/a_193_47# _1011_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X5133 VPWR _1011_/a_1059_315# _1011_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5134 _1011_/a_1017_47# _1011_/a_27_47# _1011_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X5135 _1011_/a_193_47# _1011_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X5136 _1011_/a_466_413# _1011_/a_27_47# _1011_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X5137 VGND _1011_/a_891_413# _1011_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5138 _1011_/a_381_47# _0109_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5139 VGND net97 _1011_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5140 _0726_/a_240_47# net227 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X5141 _0109_ _0726_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X5142 VGND _0219_ _0726_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5143 _0726_/a_51_297# _0355_ _0726_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X5144 _0726_/a_149_47# _0345_ _0726_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X5145 _0726_/a_240_47# _0354_ _0726_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5146 VPWR _0219_ _0726_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X5147 _0109_ _0726_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X5148 _0726_/a_149_47# _0355_ _0726_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5149 _0726_/a_245_297# _0354_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5150 VPWR _0345_ _0726_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5151 _0726_/a_512_297# net227 _0726_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5152 VPWR acc0.A\[30\] _0220_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5153 _0220_ acc0.A\[30\] _0588_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X5154 _0588_/a_113_47# net59 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5155 _0220_ net59 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5156 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5157 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5158 VPWR acc0.A\[9\] _0657_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X5159 VGND acc0.A\[9\] _0289_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X5160 _0657_/a_109_297# net67 _0289_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5161 _0289_ net67 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5162 _0511_/a_81_21# _0187_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X5163 _0511_/a_299_297# _0187_ _0511_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X5164 VPWR _0511_/a_81_21# _0156_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5165 VPWR net192 _0511_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5166 VGND _0511_/a_81_21# _0156_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5167 VGND _0179_ _0511_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X5168 _0511_/a_299_297# _0179_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5169 _0511_/a_384_47# net192 _0511_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5170 net80 clknet_1_1__leaf__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X5171 VGND clknet_1_1__leaf__0459_ net80 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X5172 net80 clknet_1_1__leaf__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5173 VPWR clknet_1_1__leaf__0459_ net80 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5174 VPWR acc0.A\[31\] _0341_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5175 _0341_ acc0.A\[31\] _0709_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X5176 _0709_/a_113_47# net60 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5177 _0341_ net60 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5178 net67 _0991_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5179 _0991_/a_891_413# _0991_/a_193_47# _0991_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X5180 _0991_/a_561_413# _0991_/a_27_47# _0991_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X5181 VPWR net77 _0991_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X5182 net67 _0991_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5183 _0991_/a_381_47# _0089_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X5184 VGND _0991_/a_634_159# _0991_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X5185 VPWR _0991_/a_891_413# _0991_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5186 _0991_/a_466_413# _0991_/a_193_47# _0991_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5187 VPWR _0991_/a_634_159# _0991_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5188 _0991_/a_634_159# _0991_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X5189 _0991_/a_634_159# _0991_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X5190 _0991_/a_975_413# _0991_/a_193_47# _0991_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X5191 VGND _0991_/a_1059_315# _0991_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X5192 _0991_/a_193_47# _0991_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X5193 _0991_/a_891_413# _0991_/a_27_47# _0991_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5194 _0991_/a_592_47# _0991_/a_193_47# _0991_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X5195 VPWR _0991_/a_1059_315# _0991_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5196 _0991_/a_1017_47# _0991_/a_27_47# _0991_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X5197 _0991_/a_193_47# _0991_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X5198 _0991_/a_466_413# _0991_/a_27_47# _0991_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X5199 VGND _0991_/a_891_413# _0991_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5200 _0991_/a_381_47# _0089_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5201 VGND net77 _0991_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5202 net114 clknet_1_1__leaf__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X5203 VGND clknet_1_1__leaf__0462_ net114 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X5204 net114 clknet_1_1__leaf__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5205 VPWR clknet_1_1__leaf__0462_ net114 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5206 VPWR A[2] input9/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5207 net9 input9/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5208 net9 input9/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5209 VGND A[2] input9/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5210 _0974_/a_222_93# _0468_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X5211 VPWR net159 _0974_/a_544_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X5212 VGND _0974_/a_79_199# _0166_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5213 _0974_/a_222_93# _0468_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0 ps=0 w=0.42 l=0.15
X5214 VGND _0486_ _0974_/a_448_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.38675 ps=3.79 w=0.65 l=0.15
X5215 _0974_/a_448_47# _0974_/a_222_93# _0974_/a_79_199# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5216 _0974_/a_79_199# _0974_/a_222_93# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0 ps=0 w=1 l=0.15
X5217 _0974_/a_544_297# _0486_ _0974_/a_79_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5218 _0974_/a_448_47# net159 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5219 VPWR _0974_/a_79_199# _0166_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5220 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5221 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5222 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5223 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5224 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X5225 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X5226 VGND _0318_ _0690_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X5227 _0690_/a_68_297# _0321_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5228 _0322_ _0690_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5229 VPWR _0318_ _0690_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X5230 _0322_ _0690_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X5231 _0690_/a_150_297# _0321_ _0690_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5232 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X5233 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X5234 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5235 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5236 VPWR _0475_ _0957_/a_304_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.135 ps=1.27 w=1 l=0.15
X5237 _0957_/a_304_297# _0472_ _0957_/a_220_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5238 VGND _0474_ _0957_/a_32_297# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X5239 _0957_/a_220_297# _0474_ _0957_/a_114_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X5240 _0957_/a_32_297# _0473_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.169 ps=1.82 w=0.65 l=0.15
X5241 _0957_/a_32_297# _0472_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5242 VPWR _0957_/a_32_297# _0476_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X5243 _0476_ _0957_/a_32_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5244 VGND _0475_ _0957_/a_32_297# VGND sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X5245 VPWR _0957_/a_32_297# _0476_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5246 _0476_ _0957_/a_32_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.1235 ps=1.03 w=0.65 l=0.15
X5247 _0476_ _0957_/a_32_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5248 _0476_ _0957_/a_32_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X5249 _0957_/a_114_297# _0473_ _0957_/a_32_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.26 ps=2.52 w=1 l=0.15
X5250 VGND _0957_/a_32_297# _0476_ VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5251 VGND _0957_/a_32_297# _0476_ VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X5252 net74 clknet_1_1__leaf__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X5253 VGND clknet_1_1__leaf__0458_ net74 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X5254 net74 clknet_1_1__leaf__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5255 VPWR clknet_1_1__leaf__0458_ net74 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5256 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5257 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5258 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5259 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5260 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X5261 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X5262 _0673_/a_103_199# _0304_ _0673_/a_253_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.39 ps=3.8 w=0.65 l=0.15
X5263 VPWR _0673_/a_103_199# _0305_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.36 ps=2.72 w=1 l=0.15
X5264 _0673_/a_337_297# _0289_ _0673_/a_253_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.33 pd=2.66 as=0.27 ps=2.54 w=1 l=0.15
X5265 _0673_/a_103_199# _0295_ _0673_/a_337_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.425 pd=2.85 as=0 ps=0 w=1 l=0.15
X5266 _0673_/a_253_297# _0287_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5267 VPWR _0304_ _0673_/a_103_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5268 VGND _0673_/a_103_199# _0305_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.234 ps=2.02 w=0.65 l=0.15
X5269 _0673_/a_253_47# _0287_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5270 _0673_/a_253_47# _0295_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5271 VGND _0289_ _0673_/a_253_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5272 VPWR input12/a_75_212# net12 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5273 input12/a_75_212# A[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5274 input12/a_75_212# A[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5275 VGND input12/a_75_212# net12 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5276 VPWR rst input34/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5277 net34 input34/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5278 net34 input34/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5279 VGND rst input34/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5280 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5281 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5282 VPWR input23/a_75_212# net23 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5283 input23/a_75_212# B[15] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5284 input23/a_75_212# B[15] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5285 VGND input23/a_75_212# net23 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5286 VPWR clknet_0__0465_ clkbuf_1_0__f__0465_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X5287 VPWR clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X5288 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5289 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5290 VPWR clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5291 VPWR clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5292 clkbuf_1_0__f__0465_/a_110_47# clknet_0__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5293 clkbuf_1_0__f__0465_/a_110_47# clknet_0__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X5294 VGND clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X5295 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5296 VGND clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5297 clkbuf_1_0__f__0465_/a_110_47# clknet_0__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5298 VGND clknet_0__0465_ clkbuf_1_0__f__0465_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5299 VGND clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5300 VPWR clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5301 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5302 VGND clknet_0__0465_ clkbuf_1_0__f__0465_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5303 VGND clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5304 VPWR clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5305 VGND clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5306 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5307 clkbuf_1_0__f__0465_/a_110_47# clknet_0__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5308 VPWR clknet_0__0465_ clkbuf_1_0__f__0465_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5309 VPWR clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5310 VPWR clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5311 VGND clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5312 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5313 VGND clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5314 VGND clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5315 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5316 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5317 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5318 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5319 VPWR clkbuf_1_0__f__0465_/a_110_47# clknet_1_0__leaf__0465_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5320 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5321 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5322 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5323 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5324 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5325 clknet_1_0__leaf__0465_ clkbuf_1_0__f__0465_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5326 _0742_/a_81_21# _0343_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X5327 _0742_/a_299_297# _0343_ _0742_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X5328 VPWR _0742_/a_81_21# _0368_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5329 VPWR _0315_ _0742_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5330 VGND _0742_/a_81_21# _0368_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5331 VGND _0366_ _0742_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X5332 _0742_/a_299_297# _0366_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5333 _0742_/a_384_47# _0315_ _0742_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5334 _0811_/a_81_21# _0346_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X5335 _0811_/a_299_297# _0346_ _0811_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X5336 VPWR _0811_/a_81_21# _0422_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5337 VPWR _0402_ _0811_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5338 VGND _0811_/a_81_21# _0422_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5339 VGND _0421_ _0811_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X5340 _0811_/a_299_297# _0421_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5341 _0811_/a_384_47# _0402_ _0811_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5342 net56 _1010_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5343 _1010_/a_891_413# _1010_/a_193_47# _1010_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X5344 _1010_/a_561_413# _1010_/a_27_47# _1010_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X5345 VPWR net96 _1010_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X5346 net56 _1010_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5347 _1010_/a_381_47# _0108_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X5348 VGND _1010_/a_634_159# _1010_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X5349 VPWR _1010_/a_891_413# _1010_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5350 _1010_/a_466_413# _1010_/a_193_47# _1010_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5351 VPWR _1010_/a_634_159# _1010_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5352 _1010_/a_634_159# _1010_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X5353 _1010_/a_634_159# _1010_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X5354 _1010_/a_975_413# _1010_/a_193_47# _1010_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X5355 VGND _1010_/a_1059_315# _1010_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X5356 _1010_/a_193_47# _1010_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X5357 _1010_/a_891_413# _1010_/a_27_47# _1010_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5358 _1010_/a_592_47# _1010_/a_193_47# _1010_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X5359 VPWR _1010_/a_1059_315# _1010_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5360 _1010_/a_1017_47# _1010_/a_27_47# _1010_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X5361 _1010_/a_193_47# _1010_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X5362 _1010_/a_466_413# _1010_/a_27_47# _1010_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X5363 VGND _1010_/a_891_413# _1010_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5364 _1010_/a_381_47# _0108_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5365 VGND net96 _1010_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5366 VPWR _0725_/a_80_21# _0355_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X5367 _0725_/a_209_297# _0353_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.65 pd=5.3 as=0 ps=0 w=1 l=0.15
X5368 _0725_/a_303_47# _0333_ _0725_/a_209_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.208 ps=1.94 w=0.65 l=0.15
X5369 _0725_/a_209_47# _0353_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5370 VGND _0725_/a_80_21# _0355_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.17225 ps=1.83 w=0.65 l=0.15
X5371 VGND _0343_ _0725_/a_80_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2145 ps=1.96 w=0.65 l=0.15
X5372 _0725_/a_80_21# _0221_ _0725_/a_303_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5373 VPWR _0333_ _0725_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5374 _0725_/a_80_21# _0343_ _0725_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0 ps=0 w=1 l=0.15
X5375 _0725_/a_209_297# _0221_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5376 VPWR net67 _0656_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X5377 _0288_ _0656_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X5378 VGND net67 _0656_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X5379 _0656_/a_59_75# acc0.A\[9\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5380 _0288_ _0656_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X5381 _0656_/a_145_75# acc0.A\[9\] _0656_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X5382 VPWR _0218_ _0587_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X5383 VGND _0587_/a_27_47# _0219_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X5384 VGND _0587_/a_27_47# _0219_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5385 _0219_ _0587_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X5386 _0219_ _0587_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5387 VGND _0218_ _0587_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X5388 VPWR _0587_/a_27_47# _0219_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5389 _0219_ _0587_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5390 _0219_ _0587_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5391 VPWR _0587_/a_27_47# _0219_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5392 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X5393 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X5394 VPWR net4 _0510_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X5395 _0510_/a_27_297# _0186_ _0510_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X5396 VGND net4 _0510_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X5397 _0187_ _0510_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5398 _0510_/a_27_297# _0186_ _0510_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X5399 _0510_/a_109_297# _0181_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5400 _0510_/a_373_47# _0181_ _0510_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5401 _0187_ _0510_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5402 _0510_/a_109_297# acc0.A\[12\] _0510_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5403 _0510_/a_109_47# acc0.A\[12\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5404 VPWR acc0.A\[5\] hold1/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5405 VGND hold1/a_285_47# hold1/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X5406 net148 hold1/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5407 VGND acc0.A\[5\] hold1/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5408 VPWR hold1/a_285_47# hold1/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X5409 hold1/a_285_47# hold1/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X5410 hold1/a_285_47# hold1/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X5411 net148 hold1/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5412 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5413 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5414 VGND acc0.A\[31\] _0708_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X5415 _0708_/a_68_297# net60 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5416 _0340_ _0708_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5417 VPWR acc0.A\[31\] _0708_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X5418 _0340_ _0708_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X5419 _0708_/a_150_297# net60 _0708_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5420 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5421 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5422 VPWR _0256_ _0639_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X5423 VGND _0256_ _0271_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X5424 _0639_/a_109_297# _0270_ _0271_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5425 _0271_ _0270_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5426 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X5427 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X5428 net66 _0990_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5429 _0990_/a_891_413# _0990_/a_193_47# _0990_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X5430 _0990_/a_561_413# _0990_/a_27_47# _0990_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X5431 VPWR net76 _0990_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X5432 net66 _0990_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5433 _0990_/a_381_47# _0088_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X5434 VGND _0990_/a_634_159# _0990_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X5435 VPWR _0990_/a_891_413# _0990_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5436 _0990_/a_466_413# _0990_/a_193_47# _0990_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5437 VPWR _0990_/a_634_159# _0990_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5438 _0990_/a_634_159# _0990_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X5439 _0990_/a_634_159# _0990_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X5440 _0990_/a_975_413# _0990_/a_193_47# _0990_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X5441 VGND _0990_/a_1059_315# _0990_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X5442 _0990_/a_193_47# _0990_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X5443 _0990_/a_891_413# _0990_/a_27_47# _0990_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5444 _0990_/a_592_47# _0990_/a_193_47# _0990_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X5445 VPWR _0990_/a_1059_315# _0990_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5446 _0990_/a_1017_47# _0990_/a_27_47# _0990_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X5447 _0990_/a_193_47# _0990_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X5448 _0990_/a_466_413# _0990_/a_27_47# _0990_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X5449 VGND _0990_/a_891_413# _0990_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5450 _0990_/a_381_47# _0088_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5451 VGND net76 _0990_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5452 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5453 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5454 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5455 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5456 net118 clknet_1_1__leaf__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X5457 VGND clknet_1_1__leaf__0463_ net118 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X5458 net118 clknet_1_1__leaf__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5459 VPWR clknet_1_1__leaf__0463_ net118 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5460 VPWR _0161_ _0973_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X5461 _0973_/a_27_297# _0487_ _0973_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X5462 VGND _0161_ _0973_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X5463 _0165_ _0973_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5464 _0973_/a_27_297# _0487_ _0973_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X5465 _0973_/a_109_297# net240 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5466 _0973_/a_373_47# net240 _0973_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5467 _0165_ _0973_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5468 _0973_/a_109_297# _0369_ _0973_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5469 _0973_/a_109_47# _0369_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5470 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5471 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5472 VPWR comp0.B\[2\] _0956_/a_304_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5473 _0956_/a_304_297# comp0.B\[1\] _0956_/a_220_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5474 VGND comp0.B\[0\] _0956_/a_32_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.4225 ps=3.9 w=0.65 l=0.15
X5475 _0956_/a_220_297# comp0.B\[0\] _0956_/a_114_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.38 ps=2.76 w=1 l=0.15
X5476 _0956_/a_32_297# comp0.B\[15\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5477 _0956_/a_32_297# comp0.B\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5478 VPWR _0956_/a_32_297# _0475_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.54 ps=5.08 w=1 l=0.15
X5479 _0475_ _0956_/a_32_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5480 VGND comp0.B\[2\] _0956_/a_32_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5481 VPWR _0956_/a_32_297# _0475_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5482 _0475_ _0956_/a_32_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X5483 _0475_ _0956_/a_32_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5484 _0475_ _0956_/a_32_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5485 _0956_/a_114_297# comp0.B\[15\] _0956_/a_32_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5486 VGND _0956_/a_32_297# _0475_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5487 VGND _0956_/a_32_297# _0475_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5488 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5489 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5490 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5491 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5492 VPWR _0283_ _0421_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5493 _0421_ _0283_ _0810_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X5494 _0810_/a_113_47# _0420_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5495 _0421_ _0420_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5496 VPWR input13/a_75_212# net13 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5497 input13/a_75_212# A[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5498 input13/a_75_212# A[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5499 VGND input13/a_75_212# net13 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5500 VPWR input24/a_75_212# net24 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5501 input24/a_75_212# B[1] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5502 input24/a_75_212# B[1] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5503 VGND input24/a_75_212# net24 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5504 VPWR clknet_0__0464_ clkbuf_1_0__f__0464_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X5505 VPWR clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X5506 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5507 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5508 VPWR clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5509 VPWR clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5510 clkbuf_1_0__f__0464_/a_110_47# clknet_0__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5511 clkbuf_1_0__f__0464_/a_110_47# clknet_0__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X5512 VGND clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X5513 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5514 VGND clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5515 clkbuf_1_0__f__0464_/a_110_47# clknet_0__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5516 VGND clknet_0__0464_ clkbuf_1_0__f__0464_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5517 VGND clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5518 VPWR clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5519 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5520 VGND clknet_0__0464_ clkbuf_1_0__f__0464_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5521 VGND clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5522 VPWR clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5523 VGND clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5524 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5525 clkbuf_1_0__f__0464_/a_110_47# clknet_0__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5526 VPWR clknet_0__0464_ clkbuf_1_0__f__0464_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5527 VPWR clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5528 VPWR clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5529 VGND clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5530 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5531 VGND clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5532 VGND clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5533 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5534 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5535 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5536 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5537 VPWR clkbuf_1_0__f__0464_/a_110_47# clknet_1_0__leaf__0464_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5538 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5539 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5540 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5541 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5542 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5543 clknet_1_0__leaf__0464_ clkbuf_1_0__f__0464_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5544 VPWR _0315_ _0741_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X5545 VGND _0315_ _0367_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X5546 _0741_/a_109_297# _0366_ _0367_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5547 _0367_ _0366_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5548 VGND _0280_ _0672_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X5549 _0672_/a_510_47# _0301_ _0672_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X5550 _0672_/a_79_21# _0303_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X5551 VPWR _0301_ _0672_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5552 _0672_/a_79_21# _0296_ _0672_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X5553 _0672_/a_297_297# _0280_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5554 _0672_/a_79_21# _0303_ _0672_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X5555 VPWR _0672_/a_79_21# _0304_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5556 VGND _0672_/a_79_21# _0304_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5557 _0672_/a_215_47# _0296_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5558 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X5559 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X5560 _0655_/a_109_93# _0286_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X5561 _0655_/a_215_53# _0283_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2226 pd=2.74 as=0 ps=0 w=0.42 l=0.15
X5562 VGND _0655_/a_109_93# _0655_/a_215_53# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5563 VGND _0280_ _0655_/a_215_53# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5564 VPWR _0280_ _0655_/a_369_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1365 ps=1.49 w=0.42 l=0.15
X5565 _0655_/a_369_297# _0283_ _0655_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X5566 _0287_ _0655_/a_215_53# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0 ps=0 w=1 l=0.15
X5567 _0655_/a_297_297# _0655_/a_109_93# _0655_/a_215_53# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5568 _0655_/a_109_93# _0286_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X5569 _0287_ _0655_/a_215_53# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X5570 VPWR _0586_/a_27_47# _0218_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5571 _0218_ _0586_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5572 VPWR control0.add _0586_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X5573 _0218_ _0586_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X5574 VGND _0586_/a_27_47# _0218_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5575 VGND control0.add _0586_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5576 _0724_/a_199_47# _0221_ _0354_ VGND sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.182 ps=1.86 w=0.65 l=0.15
X5577 _0724_/a_113_297# _0333_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.545 pd=5.09 as=0 ps=0 w=1 l=0.15
X5578 _0354_ _0353_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5579 VPWR _0221_ _0724_/a_113_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5580 _0724_/a_113_297# _0353_ _0354_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X5581 VGND _0333_ _0724_/a_199_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5582 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X5583 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X5584 control0.count\[0\] _1069_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5585 _1069_/a_891_413# _1069_/a_193_47# _1069_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X5586 _1069_/a_561_413# _1069_/a_27_47# _1069_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X5587 VPWR clknet_1_0__leaf_clk _1069_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X5588 control0.count\[0\] _1069_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5589 _1069_/a_381_47# _0167_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X5590 VGND _1069_/a_634_159# _1069_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X5591 VPWR _1069_/a_891_413# _1069_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5592 _1069_/a_466_413# _1069_/a_193_47# _1069_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5593 VPWR _1069_/a_634_159# _1069_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5594 _1069_/a_634_159# _1069_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X5595 _1069_/a_634_159# _1069_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X5596 _1069_/a_975_413# _1069_/a_193_47# _1069_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X5597 VGND _1069_/a_1059_315# _1069_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X5598 _1069_/a_193_47# _1069_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X5599 _1069_/a_891_413# _1069_/a_27_47# _1069_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5600 _1069_/a_592_47# _1069_/a_193_47# _1069_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X5601 VPWR _1069_/a_1059_315# _1069_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5602 _1069_/a_1017_47# _1069_/a_27_47# _1069_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X5603 _1069_/a_193_47# _1069_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X5604 _1069_/a_466_413# _1069_/a_27_47# _1069_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X5605 VGND _1069_/a_891_413# _1069_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5606 _1069_/a_381_47# _0167_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5607 VGND clknet_1_0__leaf_clk _1069_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5608 VPWR acc0.A\[0\] hold2/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5609 VGND hold2/a_285_47# hold2/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X5610 net149 hold2/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5611 VGND acc0.A\[0\] hold2/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5612 VPWR hold2/a_285_47# hold2/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X5613 hold2/a_285_47# hold2/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X5614 hold2/a_285_47# hold2/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X5615 net149 hold2/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5616 _0707_/a_75_199# _0338_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.38025 pd=3.77 as=0 ps=0 w=0.65 l=0.15
X5617 _0707_/a_208_47# _0334_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.25025 pd=2.07 as=0 ps=0 w=0.65 l=0.15
X5618 _0707_/a_315_47# _0333_ _0707_/a_208_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=2.34 as=0 ps=0 w=0.65 l=0.15
X5619 VGND _0335_ _0707_/a_75_199# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5620 _0707_/a_75_199# _0221_ _0707_/a_315_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5621 _0707_/a_75_199# _0338_ _0707_/a_544_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.415 ps=2.83 w=1 l=0.15
X5622 _0707_/a_544_297# _0335_ _0707_/a_201_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.655 ps=5.31 w=1 l=0.15
X5623 VPWR _0707_/a_75_199# _0339_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.285 ps=2.57 w=1 l=0.15
X5624 _0707_/a_201_297# _0334_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5625 VPWR _0333_ _0707_/a_201_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5626 _0707_/a_201_297# _0221_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5627 VGND _0707_/a_75_199# _0339_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5628 VPWR _0216_ _0569_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X5629 _0569_/a_27_297# _0195_ _0569_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X5630 VGND _0216_ _0569_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X5631 _0127_ _0569_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5632 _0569_/a_27_297# _0195_ _0569_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X5633 _0569_/a_109_297# acc0.A\[29\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5634 _0569_/a_373_47# acc0.A\[29\] _0569_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5635 _0127_ _0569_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5636 _0569_/a_109_297# net190 _0569_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5637 _0569_/a_109_47# net190 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5638 VPWR acc0.A\[4\] _0638_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X5639 VGND acc0.A\[4\] _0270_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X5640 _0638_/a_109_297# net62 _0270_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5641 _0270_ net62 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5642 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5643 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5644 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5645 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5646 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5647 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5648 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5649 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5650 _0972_/a_93_21# control0.state\[1\] _0972_/a_346_47# VGND sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.09 as=0.14625 ps=1.1 w=0.65 l=0.15
X5651 _0972_/a_93_21# _0487_ _0972_/a_250_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.185 ps=1.37 w=1 l=0.15
X5652 _0972_/a_584_47# _0487_ _0972_/a_93_21# VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.143 ps=1.09 w=0.65 l=0.15
X5653 VPWR _0972_/a_93_21# _0164_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2425 pd=1.485 as=0.33 ps=2.66 w=1 l=0.15
X5654 VGND net231 _0972_/a_584_47# VGND sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.06825 ps=0.86 w=0.65 l=0.15
X5655 _0972_/a_256_47# _0468_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0975 pd=0.95 as=0.16737 ps=1.165 w=0.65 l=0.15
X5656 _0972_/a_250_297# net231 _0972_/a_93_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X5657 VGND _0972_/a_93_21# _0164_ VGND sky130_fd_pr__nfet_01v8 ad=0.16737 pd=1.165 as=0.2145 ps=1.96 w=0.65 l=0.15
X5658 _0972_/a_250_297# _0468_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.2425 ps=1.485 w=1 l=0.15
X5659 VPWR _0471_ _0972_/a_250_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.45 as=0.165 ps=1.33 w=1 l=0.15
X5660 _0972_/a_250_297# control0.state\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.185 pd=1.37 as=0.225 ps=1.45 w=1 l=0.15
X5661 _0972_/a_346_47# _0471_ _0972_/a_256_47# VGND sky130_fd_pr__nfet_01v8 ad=0.14625 pd=1.1 as=0.0975 ps=0.95 w=0.65 l=0.15
X5662 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5663 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5664 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5665 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5666 VPWR comp0.B\[6\] _0955_/a_304_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5667 _0955_/a_304_297# comp0.B\[5\] _0955_/a_220_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5668 VGND comp0.B\[4\] _0955_/a_32_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.4225 ps=3.9 w=0.65 l=0.15
X5669 _0955_/a_220_297# comp0.B\[4\] _0955_/a_114_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.38 ps=2.76 w=1 l=0.15
X5670 _0955_/a_32_297# comp0.B\[3\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5671 _0955_/a_32_297# comp0.B\[5\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5672 VPWR _0955_/a_32_297# _0474_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.54 ps=5.08 w=1 l=0.15
X5673 _0474_ _0955_/a_32_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5674 VGND comp0.B\[6\] _0955_/a_32_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5675 VPWR _0955_/a_32_297# _0474_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5676 _0474_ _0955_/a_32_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X5677 _0474_ _0955_/a_32_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5678 _0474_ _0955_/a_32_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5679 _0955_/a_114_297# comp0.B\[3\] _0955_/a_32_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5680 VGND _0955_/a_32_297# _0474_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5681 VGND _0955_/a_32_297# _0474_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5682 VPWR _0324_ _0366_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5683 _0366_ _0324_ _0740_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X5684 _0740_/a_113_47# _0359_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5685 _0366_ _0359_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5686 VPWR input14/a_75_212# net14 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5687 input14/a_75_212# A[7] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5688 input14/a_75_212# A[7] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5689 VGND input14/a_75_212# net14 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5690 VPWR input25/a_75_212# net25 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5691 input25/a_75_212# B[2] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5692 input25/a_75_212# B[2] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5693 VGND input25/a_75_212# net25 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5694 VPWR clknet_0__0463_ clkbuf_1_0__f__0463_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X5695 VPWR clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X5696 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5697 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5698 VPWR clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5699 VPWR clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5700 clkbuf_1_0__f__0463_/a_110_47# clknet_0__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5701 clkbuf_1_0__f__0463_/a_110_47# clknet_0__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X5702 VGND clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X5703 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5704 VGND clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5705 clkbuf_1_0__f__0463_/a_110_47# clknet_0__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5706 VGND clknet_0__0463_ clkbuf_1_0__f__0463_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5707 VGND clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5708 VPWR clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5709 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5710 VGND clknet_0__0463_ clkbuf_1_0__f__0463_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5711 VGND clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5712 VPWR clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5713 VGND clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5714 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5715 clkbuf_1_0__f__0463_/a_110_47# clknet_0__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5716 VPWR clknet_0__0463_ clkbuf_1_0__f__0463_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5717 VPWR clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5718 VPWR clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5719 VGND clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5720 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5721 VGND clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5722 VGND clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5723 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5724 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5725 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5726 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5727 VPWR clkbuf_1_0__f__0463_/a_110_47# clknet_1_0__leaf__0463_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5728 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5729 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5730 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5731 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5732 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5733 clknet_1_0__leaf__0463_ clkbuf_1_0__f__0463_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5734 _0671_/a_199_47# acc0.A\[15\] _0303_ VGND sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.182 ps=1.86 w=0.65 l=0.15
X5735 _0671_/a_113_297# net42 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.545 pd=5.09 as=0 ps=0 w=1 l=0.15
X5736 _0303_ _0302_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5737 VPWR acc0.A\[15\] _0671_/a_113_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5738 _0671_/a_113_297# _0302_ _0303_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X5739 VGND net42 _0671_/a_199_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5740 VPWR clknet_1_0__leaf__0457_ _0869_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5741 _0459_ _0869_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5742 _0459_ _0869_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5743 VGND clknet_1_0__leaf__0457_ _0869_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5744 net91 clknet_1_0__leaf__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X5745 VGND clknet_1_0__leaf__0460_ net91 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X5746 net91 clknet_1_0__leaf__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5747 VPWR clknet_1_0__leaf__0460_ net91 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5748 VPWR _0334_ _0723_/a_207_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1218 ps=1.42 w=0.42 l=0.15
X5749 _0353_ _0723_/a_207_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5750 _0723_/a_297_47# _0723_/a_27_413# _0723_/a_207_413# VGND sky130_fd_pr__nfet_01v8 ad=0.1008 pd=1.32 as=0.1092 ps=1.36 w=0.42 l=0.15
X5751 _0353_ _0723_/a_207_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5752 _0723_/a_207_413# _0723_/a_27_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5753 VPWR _0335_ _0723_/a_27_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5754 VGND _0334_ _0723_/a_297_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5755 _0723_/a_27_413# _0335_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X5756 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5757 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5758 VPWR _0285_ _0654_/a_207_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1218 ps=1.42 w=0.42 l=0.15
X5759 _0286_ _0654_/a_207_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5760 _0654_/a_297_47# _0654_/a_27_413# _0654_/a_207_413# VGND sky130_fd_pr__nfet_01v8 ad=0.1008 pd=1.32 as=0.1092 ps=1.36 w=0.42 l=0.15
X5761 _0286_ _0654_/a_207_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5762 _0654_/a_207_413# _0654_/a_27_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5763 VPWR _0284_ _0654_/a_27_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5764 VGND _0285_ _0654_/a_297_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5765 _0654_/a_27_413# _0284_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X5766 VPWR net1 _0585_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X5767 _0585_/a_27_297# _0216_ _0585_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X5768 VGND net1 _0585_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X5769 _0112_ _0585_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5770 _0585_/a_27_297# _0216_ _0585_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X5771 _0585_/a_109_297# _0181_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5772 _0585_/a_373_47# _0181_ _0585_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5773 _0112_ _0585_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5774 _0585_/a_109_297# net149 _0585_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5775 _0585_/a_109_47# net149 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5776 net35 _1068_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5777 _1068_/a_891_413# _1068_/a_193_47# _1068_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X5778 _1068_/a_561_413# _1068_/a_27_47# _1068_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X5779 VPWR clknet_1_0__leaf_clk _1068_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X5780 net35 _1068_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5781 _1068_/a_381_47# _0166_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X5782 VGND _1068_/a_634_159# _1068_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X5783 VPWR _1068_/a_891_413# _1068_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5784 _1068_/a_466_413# _1068_/a_193_47# _1068_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5785 VPWR _1068_/a_634_159# _1068_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5786 _1068_/a_634_159# _1068_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X5787 _1068_/a_634_159# _1068_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X5788 _1068_/a_975_413# _1068_/a_193_47# _1068_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X5789 VGND _1068_/a_1059_315# _1068_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X5790 _1068_/a_193_47# _1068_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X5791 _1068_/a_891_413# _1068_/a_27_47# _1068_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5792 _1068_/a_592_47# _1068_/a_193_47# _1068_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X5793 VPWR _1068_/a_1059_315# _1068_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5794 _1068_/a_1017_47# _1068_/a_27_47# _1068_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X5795 _1068_/a_193_47# _1068_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X5796 _1068_/a_466_413# _1068_/a_27_47# _1068_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X5797 VGND _1068_/a_891_413# _1068_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5798 _1068_/a_381_47# _0166_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5799 VGND clknet_1_0__leaf_clk _1068_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5800 VPWR acc0.A\[21\] hold3/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5801 VGND hold3/a_285_47# hold3/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X5802 net150 hold3/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5803 VGND acc0.A\[21\] hold3/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5804 VPWR hold3/a_285_47# hold3/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X5805 hold3/a_285_47# hold3/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X5806 hold3/a_285_47# hold3/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X5807 net150 hold3/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5808 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X5809 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X5810 _0338_ _0337_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X5811 VGND _0337_ _0338_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X5812 _0338_ _0337_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5813 VPWR _0337_ _0338_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5814 _0637_/a_56_297# _0263_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.545 pd=5.09 as=0 ps=0 w=1 l=0.15
X5815 VPWR _0267_ _0637_/a_56_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5816 _0269_ _0261_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.35425 pd=3.69 as=0 ps=0 w=0.65 l=0.15
X5817 _0637_/a_139_47# _0267_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X5818 _0637_/a_311_297# _0268_ _0637_/a_56_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.31 pd=2.62 as=0 ps=0 w=1 l=0.15
X5819 _0269_ _0261_ _0637_/a_311_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0 ps=0 w=1 l=0.15
X5820 VGND _0268_ _0269_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5821 _0269_ _0263_ _0637_/a_139_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5822 VPWR _0216_ _0568_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X5823 _0568_/a_27_297# _0195_ _0568_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X5824 VGND _0216_ _0568_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X5825 _0128_ _0568_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5826 _0568_/a_27_297# _0195_ _0568_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X5827 _0568_/a_109_297# net208 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5828 _0568_/a_373_47# net208 _0568_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5829 _0128_ _0568_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5830 _0568_/a_109_297# acc0.A\[29\] _0568_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5831 _0568_/a_109_47# acc0.A\[29\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5832 VPWR control0.sh _0499_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X5833 _0178_ _0499_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X5834 VGND control0.sh _0499_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X5835 _0499_/a_59_75# _0171_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5836 _0178_ _0499_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X5837 _0499_/a_145_75# _0171_ _0499_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X5838 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X5839 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X5840 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5841 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5842 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X5843 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X5844 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X5845 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X5846 _0971_/a_81_21# _0467_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X5847 _0971_/a_299_297# _0467_ _0971_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X5848 VPWR _0971_/a_81_21# _0163_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5849 VPWR _0181_ _0971_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5850 VGND _0971_/a_81_21# _0163_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5851 VGND _0487_ _0971_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X5852 _0971_/a_299_297# _0487_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5853 _0971_/a_384_47# _0181_ _0971_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5854 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X5855 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X5856 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X5857 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X5858 VPWR comp0.B\[14\] _0954_/a_304_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5859 _0954_/a_304_297# comp0.B\[13\] _0954_/a_220_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5860 VGND comp0.B\[12\] _0954_/a_32_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.4225 ps=3.9 w=0.65 l=0.15
X5861 _0954_/a_220_297# comp0.B\[12\] _0954_/a_114_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.38 ps=2.76 w=1 l=0.15
X5862 _0954_/a_32_297# comp0.B\[11\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5863 _0954_/a_32_297# comp0.B\[13\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5864 VPWR _0954_/a_32_297# _0473_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.54 ps=5.08 w=1 l=0.15
X5865 _0473_ _0954_/a_32_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5866 VGND comp0.B\[14\] _0954_/a_32_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5867 VPWR _0954_/a_32_297# _0473_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5868 _0473_ _0954_/a_32_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X5869 _0473_ _0954_/a_32_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5870 _0473_ _0954_/a_32_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5871 _0954_/a_114_297# comp0.B\[11\] _0954_/a_32_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5872 VGND _0954_/a_32_297# _0473_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5873 VGND _0954_/a_32_297# _0473_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5874 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X5875 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X5876 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X5877 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X5878 VPWR input15/a_75_212# net15 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5879 input15/a_75_212# A[8] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5880 input15/a_75_212# A[8] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5881 VGND input15/a_75_212# net15 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5882 VPWR input26/a_75_212# net26 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X5883 input26/a_75_212# B[3] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X5884 input26/a_75_212# B[3] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X5885 VGND input26/a_75_212# net26 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X5886 VPWR clknet_0__0462_ clkbuf_1_0__f__0462_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X5887 VPWR clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X5888 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5889 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5890 VPWR clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5891 VPWR clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5892 clkbuf_1_0__f__0462_/a_110_47# clknet_0__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5893 clkbuf_1_0__f__0462_/a_110_47# clknet_0__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X5894 VGND clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X5895 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5896 VGND clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5897 clkbuf_1_0__f__0462_/a_110_47# clknet_0__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5898 VGND clknet_0__0462_ clkbuf_1_0__f__0462_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5899 VGND clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5900 VPWR clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5901 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5902 VGND clknet_0__0462_ clkbuf_1_0__f__0462_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5903 VGND clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5904 VPWR clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5905 VGND clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5906 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5907 clkbuf_1_0__f__0462_/a_110_47# clknet_0__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5908 VPWR clknet_0__0462_ clkbuf_1_0__f__0462_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5909 VPWR clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5910 VPWR clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5911 VGND clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5912 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5913 VGND clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5914 VGND clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5915 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5916 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5917 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5918 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5919 VPWR clkbuf_1_0__f__0462_/a_110_47# clknet_1_0__leaf__0462_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5920 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5921 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5922 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5923 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5924 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5925 clknet_1_0__leaf__0462_ clkbuf_1_0__f__0462_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5926 VGND acc0.A\[15\] _0670_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X5927 _0670_/a_510_47# net41 _0670_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X5928 _0670_/a_79_21# acc0.A\[14\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X5929 VPWR net41 _0670_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5930 _0670_/a_79_21# net42 _0670_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X5931 _0670_/a_297_297# acc0.A\[15\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5932 _0670_/a_79_21# acc0.A\[14\] _0670_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X5933 VPWR _0670_/a_79_21# _0302_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5934 VGND _0670_/a_79_21# _0302_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5935 _0670_/a_215_47# net42 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5936 VPWR _0799_/a_80_21# _0413_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X5937 _0799_/a_209_297# _0404_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.65 pd=5.3 as=0 ps=0 w=1 l=0.15
X5938 _0799_/a_303_47# _0298_ _0799_/a_209_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.208 ps=1.94 w=0.65 l=0.15
X5939 _0799_/a_209_47# _0404_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5940 VGND _0799_/a_80_21# _0413_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.17225 ps=1.83 w=0.65 l=0.15
X5941 VGND _0343_ _0799_/a_80_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2145 ps=1.96 w=0.65 l=0.15
X5942 _0799_/a_80_21# _0411_ _0799_/a_303_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5943 VPWR _0298_ _0799_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5944 _0799_/a_80_21# _0343_ _0799_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0 ps=0 w=1 l=0.15
X5945 _0799_/a_209_297# _0411_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5946 VPWR acc0.A\[11\] _0285_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5947 _0285_ acc0.A\[11\] _0653_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X5948 _0653_/a_113_47# net38 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5949 _0285_ net38 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5950 VGND _0347_ _0722_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X5951 _0722_/a_510_47# _0351_ _0722_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X5952 _0722_/a_79_21# _0352_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X5953 VPWR _0351_ _0722_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5954 _0722_/a_79_21# _0349_ _0722_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X5955 _0722_/a_297_297# _0347_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5956 _0722_/a_79_21# _0352_ _0722_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X5957 VPWR _0722_/a_79_21# _0110_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X5958 VGND _0722_/a_79_21# _0110_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5959 _0722_/a_215_47# _0349_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5960 VPWR net23 _0584_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X5961 _0584_/a_27_297# _0216_ _0584_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X5962 VGND net23 _0584_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X5963 _0113_ _0584_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5964 _0584_/a_27_297# _0216_ _0584_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X5965 _0584_/a_109_297# _0181_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5966 _0584_/a_373_47# _0181_ _0584_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5967 _0113_ _0584_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5968 _0584_/a_109_297# net157 _0584_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X5969 _0584_/a_109_47# net157 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X5970 control0.add _1067_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X5971 _1067_/a_891_413# _1067_/a_193_47# _1067_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X5972 _1067_/a_561_413# _1067_/a_27_47# _1067_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X5973 VPWR clknet_1_1__leaf_clk _1067_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X5974 control0.add _1067_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5975 _1067_/a_381_47# _0165_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X5976 VGND _1067_/a_634_159# _1067_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X5977 VPWR _1067_/a_891_413# _1067_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X5978 _1067_/a_466_413# _1067_/a_193_47# _1067_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5979 VPWR _1067_/a_634_159# _1067_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5980 _1067_/a_634_159# _1067_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X5981 _1067_/a_634_159# _1067_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X5982 _1067_/a_975_413# _1067_/a_193_47# _1067_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X5983 VGND _1067_/a_1059_315# _1067_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X5984 _1067_/a_193_47# _1067_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X5985 _1067_/a_891_413# _1067_/a_27_47# _1067_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5986 _1067_/a_592_47# _1067_/a_193_47# _1067_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X5987 VPWR _1067_/a_1059_315# _1067_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5988 _1067_/a_1017_47# _1067_/a_27_47# _1067_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X5989 _1067_/a_193_47# _1067_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X5990 _1067_/a_466_413# _1067_/a_27_47# _1067_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X5991 VGND _1067_/a_891_413# _1067_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X5992 _1067_/a_381_47# _0165_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X5993 VGND clknet_1_1__leaf_clk _1067_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5994 VPWR _0120_ hold4/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5995 VGND hold4/a_285_47# hold4/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X5996 net151 hold4/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X5997 VGND _0120_ hold4/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X5998 VPWR hold4/a_285_47# hold4/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X5999 hold4/a_285_47# hold4/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X6000 hold4/a_285_47# hold4/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X6001 net151 hold4/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6002 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6003 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6004 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6005 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6006 VPWR net61 _0636_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6007 _0268_ _0636_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X6008 VGND net61 _0636_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6009 _0636_/a_59_75# acc0.A\[3\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6010 _0268_ _0636_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X6011 _0636_/a_145_75# acc0.A\[3\] _0636_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X6012 VPWR _0336_ _0705_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6013 _0337_ _0705_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X6014 VGND _0336_ _0705_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6015 _0705_/a_59_75# _0220_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6016 _0337_ _0705_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X6017 _0705_/a_145_75# _0220_ _0705_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X6018 _0498_/a_240_47# net7 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X6019 _0159_ _0498_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X6020 VGND _0172_ _0498_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6021 _0498_/a_51_297# net247 _0498_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X6022 _0498_/a_149_47# _0177_ _0498_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X6023 _0498_/a_240_47# _0174_ _0498_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6024 VPWR _0172_ _0498_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X6025 _0159_ _0498_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X6026 _0498_/a_149_47# net247 _0498_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6027 _0498_/a_245_297# _0174_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6028 VPWR _0177_ _0498_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6029 _0498_/a_512_297# net7 _0498_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6030 VPWR _0216_ _0567_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X6031 _0567_/a_27_297# _0195_ _0567_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X6032 VGND _0216_ _0567_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X6033 _0129_ _0567_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6034 _0567_/a_27_297# _0195_ _0567_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X6035 _0567_/a_109_297# net162 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6036 _0567_/a_373_47# net162 _0567_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6037 _0129_ _0567_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6038 _0567_/a_109_297# acc0.A\[30\] _0567_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6039 _0567_/a_109_47# acc0.A\[30\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6040 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6041 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6042 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6043 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6044 net129 clknet_1_1__leaf__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X6045 VGND clknet_1_1__leaf__0464_ net129 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6046 net129 clknet_1_1__leaf__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6047 VPWR clknet_1_1__leaf__0464_ net129 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6048 net143 clknet_1_1__leaf__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X6049 VGND clknet_1_1__leaf__0465_ net143 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6050 net143 clknet_1_1__leaf__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6051 VPWR clknet_1_1__leaf__0465_ net143 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6052 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6053 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6054 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6055 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6056 VGND acc0.A\[7\] _0619_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6057 _0619_/a_68_297# net65 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6058 _0251_ _0619_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6059 VPWR acc0.A\[7\] _0619_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X6060 _0251_ _0619_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X6061 _0619_/a_150_297# net65 _0619_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6062 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6063 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6064 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6065 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6066 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X6067 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X6068 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X6069 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X6070 VGND _0484_ _0970_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.06825 ps=0.86 w=0.65 l=0.15
X6071 VGND _0487_ _0162_ VGND sky130_fd_pr__nfet_01v8 ad=0.26 pd=2.1 as=0.08775 ps=0.92 w=0.65 l=0.15
X6072 _0162_ _0485_ _0970_/a_114_47# VGND sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.08937 ps=0.925 w=0.65 l=0.15
X6073 _0970_/a_114_47# _0484_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08937 pd=0.925 as=0.18525 ps=1.87 w=0.65 l=0.15
X6074 _0970_/a_27_297# _0487_ _0162_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0.135 ps=1.27 w=1 l=0.15
X6075 _0970_/a_27_297# _0485_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X6076 _0162_ _0487_ _0970_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6077 VPWR _0484_ _0970_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.28 ps=2.56 w=1 l=0.15
X6078 _0970_/a_27_297# _0484_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6079 VPWR _0485_ _0970_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14 ps=1.28 w=1 l=0.15
X6080 _0970_/a_285_47# _0485_ _0162_ VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.091 ps=0.93 w=0.65 l=0.15
X6081 _0162_ _0487_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X6082 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X6083 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X6084 net110 clknet_1_0__leaf__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X6085 VGND clknet_1_0__leaf__0462_ net110 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6086 net110 clknet_1_0__leaf__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6087 VPWR clknet_1_0__leaf__0462_ net110 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6088 net124 clknet_1_0__leaf__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X6089 VGND clknet_1_0__leaf__0463_ net124 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6090 net124 clknet_1_0__leaf__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6091 VPWR clknet_1_0__leaf__0463_ net124 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6092 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6093 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6094 VPWR comp0.B\[10\] _0953_/a_304_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6095 _0953_/a_304_297# comp0.B\[9\] _0953_/a_220_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6096 VGND comp0.B\[8\] _0953_/a_32_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.4225 ps=3.9 w=0.65 l=0.15
X6097 _0953_/a_220_297# comp0.B\[8\] _0953_/a_114_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.38 ps=2.76 w=1 l=0.15
X6098 _0953_/a_32_297# comp0.B\[7\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6099 _0953_/a_32_297# comp0.B\[9\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6100 VPWR _0953_/a_32_297# _0472_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.54 ps=5.08 w=1 l=0.15
X6101 _0472_ _0953_/a_32_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6102 VGND comp0.B\[10\] _0953_/a_32_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6103 VPWR _0953_/a_32_297# _0472_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6104 _0472_ _0953_/a_32_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X6105 _0472_ _0953_/a_32_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6106 _0472_ _0953_/a_32_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6107 _0953_/a_114_297# comp0.B\[7\] _0953_/a_32_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X6108 VGND _0953_/a_32_297# _0472_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6109 VGND _0953_/a_32_297# _0472_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6110 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6111 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6112 VPWR input16/a_75_212# net16 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X6113 input16/a_75_212# A[9] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X6114 input16/a_75_212# A[9] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X6115 VGND input16/a_75_212# net16 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X6116 VPWR input27/a_75_212# net27 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X6117 input27/a_75_212# B[4] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X6118 input27/a_75_212# B[4] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X6119 VGND input27/a_75_212# net27 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X6120 VPWR clknet_0__0461_ clkbuf_1_0__f__0461_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X6121 VPWR clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X6122 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6123 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6124 VPWR clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6125 VPWR clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6126 clkbuf_1_0__f__0461_/a_110_47# clknet_0__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6127 clkbuf_1_0__f__0461_/a_110_47# clknet_0__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X6128 VGND clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X6129 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6130 VGND clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6131 clkbuf_1_0__f__0461_/a_110_47# clknet_0__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6132 VGND clknet_0__0461_ clkbuf_1_0__f__0461_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6133 VGND clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6134 VPWR clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6135 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6136 VGND clknet_0__0461_ clkbuf_1_0__f__0461_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6137 VGND clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6138 VPWR clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6139 VGND clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6140 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6141 clkbuf_1_0__f__0461_/a_110_47# clknet_0__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6142 VPWR clknet_0__0461_ clkbuf_1_0__f__0461_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6143 VPWR clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6144 VPWR clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6145 VGND clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6146 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6147 VGND clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6148 VGND clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6149 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6150 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6151 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6152 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6153 VPWR clkbuf_1_0__f__0461_/a_110_47# clknet_1_0__leaf__0461_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6154 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6155 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6156 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6157 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6158 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6159 clknet_1_0__leaf__0461_ clkbuf_1_0__f__0461_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6160 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X6161 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X6162 _0798_/a_199_47# _0298_ _0412_ VGND sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.182 ps=1.86 w=0.65 l=0.15
X6163 _0798_/a_113_297# _0404_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.545 pd=5.09 as=0 ps=0 w=1 l=0.15
X6164 _0412_ _0411_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6165 VPWR _0298_ _0798_/a_113_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6166 _0798_/a_113_297# _0411_ _0412_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X6167 VGND _0404_ _0798_/a_199_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6168 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6169 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6170 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6171 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6172 VPWR _0208_ _0721_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X6173 VGND _0721_/a_27_47# _0352_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X6174 VGND _0721_/a_27_47# _0352_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6175 _0352_ _0721_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X6176 _0352_ _0721_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6177 VGND _0208_ _0721_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X6178 VPWR _0721_/a_27_47# _0352_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6179 _0352_ _0721_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6180 _0352_ _0721_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6181 VPWR _0721_/a_27_47# _0352_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6182 VPWR _0183_ _0583_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X6183 _0583_/a_27_297# _0217_ _0583_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X6184 VGND _0183_ _0583_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X6185 _0114_ _0583_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6186 _0583_/a_27_297# _0217_ _0583_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X6187 _0583_/a_109_297# acc0.A\[16\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6188 _0583_/a_373_47# acc0.A\[16\] _0583_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6189 _0114_ _0583_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6190 _0583_/a_109_297# net165 _0583_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6191 _0583_/a_109_47# net165 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6192 VPWR acc0.A\[11\] _0652_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X6193 VGND acc0.A\[11\] _0284_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6194 _0652_/a_109_297# net38 _0284_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X6195 _0284_ net38 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6196 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6197 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6198 control0.sh _1066_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6199 _1066_/a_891_413# _1066_/a_193_47# _1066_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X6200 _1066_/a_561_413# _1066_/a_27_47# _1066_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X6201 VPWR clknet_1_1__leaf_clk _1066_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X6202 control0.sh _1066_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6203 _1066_/a_381_47# net232 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X6204 VGND _1066_/a_634_159# _1066_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X6205 VPWR _1066_/a_891_413# _1066_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6206 _1066_/a_466_413# _1066_/a_193_47# _1066_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6207 VPWR _1066_/a_634_159# _1066_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6208 _1066_/a_634_159# _1066_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X6209 _1066_/a_634_159# _1066_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X6210 _1066_/a_975_413# _1066_/a_193_47# _1066_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X6211 VGND _1066_/a_1059_315# _1066_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X6212 _1066_/a_193_47# _1066_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X6213 _1066_/a_891_413# _1066_/a_27_47# _1066_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6214 _1066_/a_592_47# _1066_/a_193_47# _1066_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X6215 VPWR _1066_/a_1059_315# _1066_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6216 _1066_/a_1017_47# _1066_/a_27_47# _1066_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X6217 _1066_/a_193_47# _1066_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X6218 _1066_/a_466_413# _1066_/a_27_47# _1066_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X6219 VGND _1066_/a_891_413# _1066_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6220 _1066_/a_381_47# net232 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6221 VGND clknet_1_1__leaf_clk _1066_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6222 VPWR comp0.B\[10\] hold5/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6223 VGND hold5/a_285_47# hold5/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X6224 net152 hold5/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6225 VGND comp0.B\[10\] hold5/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6226 VPWR hold5/a_285_47# hold5/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X6227 hold5/a_285_47# hold5/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X6228 hold5/a_285_47# hold5/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X6229 net152 hold5/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6230 VPWR _0182_ _0566_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X6231 VGND _0566_/a_27_47# _0216_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X6232 VGND _0566_/a_27_47# _0216_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6233 _0216_ _0566_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X6234 _0216_ _0566_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6235 VGND _0182_ _0566_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X6236 VPWR _0566_/a_27_47# _0216_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6237 _0216_ _0566_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6238 _0216_ _0566_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6239 VPWR _0566_/a_27_47# _0216_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6240 _0267_ _0265_ _0635_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.348 pd=2.78 as=0.21 ps=2.42 w=1 l=0.15
X6241 VPWR _0266_ _0267_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.7 l=0.15
X6242 _0635_/a_27_47# _0265_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X6243 _0267_ _0266_ _0635_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6244 _0635_/a_109_297# _0264_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6245 VGND _0264_ _0635_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6246 VGND acc0.A\[30\] _0704_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6247 _0704_/a_68_297# net59 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6248 _0336_ _0704_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6249 VPWR acc0.A\[30\] _0704_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X6250 _0336_ _0704_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X6251 _0704_/a_150_297# net59 _0704_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6252 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6253 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6254 VGND acc0.A\[15\] _0497_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6255 _0497_/a_68_297# _0176_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6256 _0177_ _0497_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6257 VPWR acc0.A\[15\] _0497_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X6258 _0177_ _0497_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X6259 _0497_/a_150_297# _0176_ _0497_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6260 acc0.A\[3\] _1049_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6261 _1049_/a_891_413# _1049_/a_193_47# _1049_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X6262 _1049_/a_561_413# _1049_/a_27_47# _1049_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X6263 VPWR net135 _1049_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X6264 acc0.A\[3\] _1049_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6265 _1049_/a_381_47# _0147_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X6266 VGND _1049_/a_634_159# _1049_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X6267 VPWR _1049_/a_891_413# _1049_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6268 _1049_/a_466_413# _1049_/a_193_47# _1049_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6269 VPWR _1049_/a_634_159# _1049_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6270 _1049_/a_634_159# _1049_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X6271 _1049_/a_634_159# _1049_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X6272 _1049_/a_975_413# _1049_/a_193_47# _1049_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X6273 VGND _1049_/a_1059_315# _1049_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X6274 _1049_/a_193_47# _1049_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X6275 _1049_/a_891_413# _1049_/a_27_47# _1049_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6276 _1049_/a_592_47# _1049_/a_193_47# _1049_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X6277 VPWR _1049_/a_1059_315# _1049_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6278 _1049_/a_1017_47# _1049_/a_27_47# _1049_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X6279 _1049_/a_193_47# _1049_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X6280 _1049_/a_466_413# _1049_/a_27_47# _1049_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X6281 VGND _1049_/a_891_413# _1049_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6282 _1049_/a_381_47# _0147_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6283 VGND net135 _1049_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6284 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X6285 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X6286 VGND _0222_ _0618_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X6287 _0618_/a_510_47# _0232_ _0618_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X6288 _0618_/a_79_21# _0249_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X6289 VPWR _0232_ _0618_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6290 _0618_/a_79_21# _0223_ _0618_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X6291 _0618_/a_297_297# _0222_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6292 _0618_/a_79_21# _0249_ _0618_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X6293 VPWR _0618_/a_79_21# _0250_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X6294 VGND _0618_/a_79_21# _0250_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6295 _0618_/a_215_47# _0223_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6296 VGND net171 _0549_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6297 _0549_/a_68_297# _0176_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6298 _0207_ _0549_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6299 VPWR net171 _0549_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X6300 _0207_ _0549_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X6301 _0549_/a_150_297# _0176_ _0549_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6302 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6303 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6304 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6305 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6306 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6307 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6308 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X6309 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X6310 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X6311 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X6312 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6313 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6314 _0471_ control0.state\[0\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X6315 VGND control0.state\[0\] _0471_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6316 _0471_ control0.state\[0\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6317 VPWR control0.state\[0\] _0471_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6318 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6319 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6320 net102 clknet_1_1__leaf__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X6321 VGND clknet_1_1__leaf__0461_ net102 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6322 net102 clknet_1_1__leaf__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6323 VPWR clknet_1_1__leaf__0461_ net102 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6324 VPWR input17/a_75_212# net17 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X6325 input17/a_75_212# B[0] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X6326 input17/a_75_212# B[0] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X6327 VGND input17/a_75_212# net17 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X6328 VPWR input28/a_75_212# net28 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X6329 input28/a_75_212# B[5] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X6330 input28/a_75_212# B[5] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X6331 VGND input28/a_75_212# net28 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X6332 VPWR clknet_0__0460_ clkbuf_1_0__f__0460_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X6333 VPWR clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X6334 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6335 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6336 VPWR clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6337 VPWR clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6338 clkbuf_1_0__f__0460_/a_110_47# clknet_0__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6339 clkbuf_1_0__f__0460_/a_110_47# clknet_0__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X6340 VGND clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X6341 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6342 VGND clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6343 clkbuf_1_0__f__0460_/a_110_47# clknet_0__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6344 VGND clknet_0__0460_ clkbuf_1_0__f__0460_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6345 VGND clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6346 VPWR clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6347 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6348 VGND clknet_0__0460_ clkbuf_1_0__f__0460_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6349 VGND clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6350 VPWR clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6351 VGND clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6352 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6353 clkbuf_1_0__f__0460_/a_110_47# clknet_0__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6354 VPWR clknet_0__0460_ clkbuf_1_0__f__0460_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6355 VPWR clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6356 VPWR clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6357 VGND clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6358 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6359 VGND clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6360 VGND clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6361 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6362 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6363 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6364 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6365 VPWR clkbuf_1_0__f__0460_/a_110_47# clknet_1_0__leaf__0460_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6366 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6367 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6368 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6369 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6370 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6371 clknet_1_0__leaf__0460_ clkbuf_1_0__f__0460_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6372 VPWR clknet_1_1__leaf__0457_ _0935_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X6373 _0465_ _0935_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X6374 _0465_ _0935_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X6375 VGND clknet_1_1__leaf__0457_ _0935_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X6376 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6377 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6378 VPWR _0299_ _0797_/a_207_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1218 ps=1.42 w=0.42 l=0.15
X6379 _0411_ _0797_/a_207_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6380 _0797_/a_297_47# _0797_/a_27_413# _0797_/a_207_413# VGND sky130_fd_pr__nfet_01v8 ad=0.1008 pd=1.32 as=0.1092 ps=1.36 w=0.42 l=0.15
X6381 _0411_ _0797_/a_207_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6382 _0797_/a_207_413# _0797_/a_27_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6383 VPWR _0297_ _0797_/a_27_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6384 VGND _0299_ _0797_/a_297_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6385 _0797_/a_27_413# _0297_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X6386 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6387 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6388 VGND _0350_ _0720_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6389 _0720_/a_68_297# net239 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6390 _0351_ _0720_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6391 VPWR _0350_ _0720_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X6392 _0351_ _0720_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X6393 _0720_/a_150_297# net239 _0720_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6394 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6395 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6396 VPWR _0281_ _0283_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6397 _0283_ _0281_ _0651_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X6398 _0651_/a_113_47# _0282_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6399 _0283_ _0282_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6400 VPWR _0183_ _0582_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X6401 _0582_/a_27_297# _0217_ _0582_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X6402 VGND _0183_ _0582_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X6403 _0115_ _0582_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6404 _0582_/a_27_297# _0217_ _0582_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X6405 _0582_/a_109_297# net219 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6406 _0582_/a_373_47# net219 _0582_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6407 _0115_ _0582_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6408 _0582_/a_109_297# net221 _0582_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6409 _0582_/a_109_47# net221 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6410 net83 clknet_1_1__leaf__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X6411 VGND clknet_1_1__leaf__0459_ net83 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6412 net83 clknet_1_1__leaf__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6413 VPWR clknet_1_1__leaf__0459_ net83 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6414 control0.reset _1065_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6415 _1065_/a_891_413# _1065_/a_193_47# _1065_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X6416 _1065_/a_561_413# _1065_/a_27_47# _1065_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X6417 VPWR clknet_1_1__leaf_clk _1065_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X6418 control0.reset _1065_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6419 _1065_/a_381_47# _0163_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X6420 VGND _1065_/a_634_159# _1065_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X6421 VPWR _1065_/a_891_413# _1065_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6422 _1065_/a_466_413# _1065_/a_193_47# _1065_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6423 VPWR _1065_/a_634_159# _1065_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6424 _1065_/a_634_159# _1065_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X6425 _1065_/a_634_159# _1065_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X6426 _1065_/a_975_413# _1065_/a_193_47# _1065_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X6427 VGND _1065_/a_1059_315# _1065_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X6428 _1065_/a_193_47# _1065_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X6429 _1065_/a_891_413# _1065_/a_27_47# _1065_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6430 _1065_/a_592_47# _1065_/a_193_47# _1065_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X6431 VPWR _1065_/a_1059_315# _1065_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6432 _1065_/a_1017_47# _1065_/a_27_47# _1065_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X6433 _1065_/a_193_47# _1065_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X6434 _1065_/a_466_413# _1065_/a_27_47# _1065_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X6435 VGND _1065_/a_891_413# _1065_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6436 _1065_/a_381_47# _0163_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6437 VGND clknet_1_1__leaf_clk _1065_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6438 VGND _0219_ _0849_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X6439 _0849_/a_510_47# _0451_ _0849_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X6440 _0849_/a_79_21# _0399_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X6441 VPWR _0451_ _0849_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6442 _0849_/a_79_21# net222 _0849_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X6443 _0849_/a_297_297# _0219_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6444 _0849_/a_79_21# _0399_ _0849_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X6445 VPWR _0849_/a_79_21# _0082_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X6446 VGND _0849_/a_79_21# _0082_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6447 _0849_/a_215_47# net222 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6448 VPWR _0139_ hold6/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6449 VGND hold6/a_285_47# hold6/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X6450 net153 hold6/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6451 VGND _0139_ hold6/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6452 VPWR hold6/a_285_47# hold6/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X6453 hold6/a_285_47# hold6/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X6454 hold6/a_285_47# hold6/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X6455 net153 hold6/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6456 VPWR acc0.A\[29\] _0703_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X6457 VGND acc0.A\[29\] _0335_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6458 _0703_/a_109_297# net57 _0335_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X6459 _0335_ net57 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6460 VPWR _0175_ _0496_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X6461 VPWR _0496_/a_27_47# _0176_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X6462 VGND _0175_ _0496_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X6463 _0176_ _0496_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X6464 _0176_ _0496_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X6465 VGND _0496_/a_27_47# _0176_ VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X6466 _0565_/a_240_47# net17 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X6467 _0130_ _0565_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X6468 VGND _0208_ _0565_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6469 _0565_/a_51_297# net201 _0565_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X6470 _0565_/a_149_47# _0215_ _0565_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X6471 _0565_/a_240_47# _0173_ _0565_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6472 VPWR _0208_ _0565_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X6473 _0130_ _0565_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X6474 _0565_/a_149_47# net201 _0565_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6475 _0565_/a_245_297# _0173_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6476 VPWR _0215_ _0565_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6477 _0565_/a_512_297# net17 _0565_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6478 VPWR acc0.A\[1\] _0266_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6479 _0266_ acc0.A\[1\] _0634_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X6480 _0634_/a_113_47# net47 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6481 _0266_ net47 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6482 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6483 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6484 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6485 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6486 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6487 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6488 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6489 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6490 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X6491 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X6492 acc0.A\[2\] _1048_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6493 _1048_/a_891_413# _1048_/a_193_47# _1048_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X6494 _1048_/a_561_413# _1048_/a_27_47# _1048_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X6495 VPWR net134 _1048_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X6496 acc0.A\[2\] _1048_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6497 _1048_/a_381_47# _0146_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X6498 VGND _1048_/a_634_159# _1048_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X6499 VPWR _1048_/a_891_413# _1048_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6500 _1048_/a_466_413# _1048_/a_193_47# _1048_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6501 VPWR _1048_/a_634_159# _1048_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6502 _1048_/a_634_159# _1048_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X6503 _1048_/a_634_159# _1048_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X6504 _1048_/a_975_413# _1048_/a_193_47# _1048_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X6505 VGND _1048_/a_1059_315# _1048_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X6506 _1048_/a_193_47# _1048_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X6507 _1048_/a_891_413# _1048_/a_27_47# _1048_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6508 _1048_/a_592_47# _1048_/a_193_47# _1048_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X6509 VPWR _1048_/a_1059_315# _1048_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6510 _1048_/a_1017_47# _1048_/a_27_47# _1048_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X6511 _1048_/a_193_47# _1048_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X6512 _1048_/a_466_413# _1048_/a_27_47# _1048_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X6513 VGND _1048_/a_891_413# _1048_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6514 _1048_/a_381_47# _0146_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6515 VGND net134 _1048_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6516 VPWR clknet_0_clk clkbuf_1_1__f_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X6517 VPWR clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X6518 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6519 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6520 VPWR clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6521 VPWR clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6522 clkbuf_1_1__f_clk/a_110_47# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6523 clkbuf_1_1__f_clk/a_110_47# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X6524 VGND clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X6525 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6526 VGND clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6527 clkbuf_1_1__f_clk/a_110_47# clknet_0_clk VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6528 VGND clknet_0_clk clkbuf_1_1__f_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6529 VGND clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6530 VPWR clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6531 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6532 VGND clknet_0_clk clkbuf_1_1__f_clk/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6533 VGND clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6534 VPWR clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6535 VGND clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6536 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6537 clkbuf_1_1__f_clk/a_110_47# clknet_0_clk VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6538 VPWR clknet_0_clk clkbuf_1_1__f_clk/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6539 VPWR clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6540 VPWR clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6541 VGND clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6542 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6543 VGND clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6544 VGND clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6545 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6546 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6547 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6548 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6549 VPWR clkbuf_1_1__f_clk/a_110_47# clknet_1_1__leaf_clk VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6550 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6551 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6552 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6553 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6554 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6555 clknet_1_1__leaf_clk clkbuf_1_1__f_clk/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6556 _0548_/a_240_47# net31 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X6557 _0138_ _0548_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X6558 VGND _0172_ _0548_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6559 _0548_/a_51_297# net173 _0548_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X6560 _0548_/a_149_47# _0206_ _0548_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X6561 _0548_/a_240_47# _0174_ _0548_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6562 VPWR _0172_ _0548_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X6563 _0138_ _0548_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X6564 _0548_/a_149_47# net173 _0548_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6565 _0548_/a_245_297# _0174_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6566 VPWR _0206_ _0548_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6567 _0548_/a_512_297# net31 _0548_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6568 VGND _0238_ _0617_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6569 _0617_/a_68_297# _0248_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6570 _0249_ _0617_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6571 VPWR _0238_ _0617_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X6572 _0249_ _0617_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X6573 _0617_/a_150_297# _0248_ _0617_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6574 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X6575 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X6576 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6577 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6578 net69 clknet_1_0__leaf__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X6579 VGND clknet_1_0__leaf__0458_ net69 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6580 net69 clknet_1_0__leaf__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6581 VPWR clknet_1_0__leaf__0458_ net69 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6582 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6583 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6584 _0951_/a_109_93# control0.state\[1\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.10785 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6585 _0470_ _0951_/a_209_311# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14222 ps=1.335 w=1 l=0.15
X6586 _0951_/a_109_93# control0.state\[1\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1087 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X6587 _0951_/a_296_53# _0951_/a_109_93# _0951_/a_209_311# VGND sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.10783 ps=1.36 w=0.42 l=0.15
X6588 VPWR comp0.B\[0\] _0951_/a_209_311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14222 pd=1.335 as=0.07438 ps=0.815 w=0.42 l=0.15
X6589 _0951_/a_368_53# _0161_ _0951_/a_296_53# VGND sky130_fd_pr__nfet_01v8 ad=0.05355 pd=0.675 as=0.0441 ps=0.63 w=0.42 l=0.15
X6590 _0470_ _0951_/a_209_311# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.12228 ps=1.08 w=0.65 l=0.15
X6591 _0951_/a_209_311# _0161_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07438 pd=0.815 as=0.0567 ps=0.69 w=0.42 l=0.15
X6592 VPWR _0951_/a_109_93# _0951_/a_209_311# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X6593 VGND comp0.B\[0\] _0951_/a_368_53# VGND sky130_fd_pr__nfet_01v8 ad=0.12228 pd=1.08 as=0.05355 ps=0.675 w=0.42 l=0.15
X6594 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X6595 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X6596 VPWR input18/a_75_212# net18 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X6597 input18/a_75_212# B[10] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X6598 input18/a_75_212# B[10] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X6599 VGND input18/a_75_212# net18 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X6600 VPWR input29/a_75_212# net29 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X6601 input29/a_75_212# B[6] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X6602 input29/a_75_212# B[6] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X6603 VGND input29/a_75_212# net29 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X6604 VGND _0369_ _0796_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X6605 _0796_/a_510_47# _0410_ _0796_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X6606 _0796_/a_79_21# _0399_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X6607 VPWR _0410_ _0796_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6608 _0796_/a_79_21# net238 _0796_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X6609 _0796_/a_297_297# _0369_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6610 _0796_/a_79_21# _0399_ _0796_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X6611 VPWR _0796_/a_79_21# _0094_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X6612 VGND _0796_/a_79_21# _0094_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6613 _0796_/a_215_47# net238 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6614 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6615 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6616 VPWR _0183_ _0581_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X6617 _0581_/a_27_297# _0217_ _0581_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X6618 VGND _0183_ _0581_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X6619 _0116_ _0581_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6620 _0581_/a_27_297# _0217_ _0581_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X6621 _0581_/a_109_297# net206 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6622 _0581_/a_373_47# net206 _0581_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6623 _0116_ _0581_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6624 _0581_/a_109_297# net219 _0581_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6625 _0581_/a_109_47# net219 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6626 VGND acc0.A\[10\] _0650_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6627 _0650_/a_68_297# net37 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6628 _0282_ _0650_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6629 VPWR acc0.A\[10\] _0650_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X6630 _0282_ _0650_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X6631 _0650_/a_150_297# net37 _0650_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6632 control0.state\[2\] _1064_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6633 _1064_/a_891_413# _1064_/a_193_47# _1064_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X6634 _1064_/a_561_413# _1064_/a_27_47# _1064_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X6635 VPWR clknet_1_0__leaf_clk _1064_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X6636 control0.state\[2\] _1064_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6637 _1064_/a_381_47# _0162_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X6638 VGND _1064_/a_634_159# _1064_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X6639 VPWR _1064_/a_891_413# _1064_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6640 _1064_/a_466_413# _1064_/a_193_47# _1064_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6641 VPWR _1064_/a_634_159# _1064_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6642 _1064_/a_634_159# _1064_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X6643 _1064_/a_634_159# _1064_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X6644 _1064_/a_975_413# _1064_/a_193_47# _1064_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X6645 VGND _1064_/a_1059_315# _1064_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X6646 _1064_/a_193_47# _1064_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X6647 _1064_/a_891_413# _1064_/a_27_47# _1064_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6648 _1064_/a_592_47# _1064_/a_193_47# _1064_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X6649 VPWR _1064_/a_1059_315# _1064_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6650 _1064_/a_1017_47# _1064_/a_27_47# _1064_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X6651 _1064_/a_193_47# _1064_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X6652 _1064_/a_466_413# _1064_/a_27_47# _1064_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X6653 VGND _1064_/a_891_413# _1064_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6654 _1064_/a_381_47# _0162_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6655 VGND clknet_1_0__leaf_clk _1064_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6656 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6657 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6658 net140 clknet_1_0__leaf__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X6659 VGND clknet_1_0__leaf__0465_ net140 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6660 net140 clknet_1_0__leaf__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6661 VPWR clknet_1_0__leaf__0465_ net140 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6662 _0451_ _0450_ _0848_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.348 pd=2.78 as=0.21 ps=2.42 w=1 l=0.15
X6663 VPWR _0350_ _0451_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.7 l=0.15
X6664 _0848_/a_27_47# _0450_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X6665 _0451_ _0350_ _0848_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6666 _0848_/a_109_297# _0446_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6667 VGND _0446_ _0848_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6668 VGND _0347_ _0779_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X6669 _0779_/a_510_47# _0396_ _0779_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X6670 _0779_/a_79_21# _0352_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X6671 VPWR _0396_ _0779_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6672 _0779_/a_79_21# _0395_ _0779_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X6673 _0779_/a_297_297# _0347_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6674 _0779_/a_79_21# _0352_ _0779_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X6675 VPWR _0779_/a_79_21# _0097_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X6676 VGND _0779_/a_79_21# _0097_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6677 _0779_/a_215_47# _0395_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6678 VPWR acc0.A\[4\] hold7/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6679 VGND hold7/a_285_47# hold7/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X6680 net154 hold7/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6681 VGND acc0.A\[4\] hold7/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6682 VPWR hold7/a_285_47# hold7/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X6683 hold7/a_285_47# hold7/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X6684 hold7/a_285_47# hold7/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X6685 net154 hold7/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6686 VPWR acc0.A\[29\] _0334_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6687 _0334_ acc0.A\[29\] _0702_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X6688 _0702_/a_113_47# net57 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6689 _0334_ net57 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6690 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6691 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6692 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6693 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6694 VPWR acc0.A\[1\] _0633_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X6695 VGND acc0.A\[1\] _0265_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6696 _0633_/a_109_297# net47 _0265_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X6697 _0265_ net47 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6698 VGND control0.reset _0495_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6699 _0495_/a_68_297# control0.sh VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6700 _0175_ _0495_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6701 VPWR control0.reset _0495_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X6702 _0175_ _0495_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X6703 _0495_/a_150_297# control0.sh _0495_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6704 VGND comp0.B\[0\] _0564_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6705 _0564_/a_68_297# _0175_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6706 _0215_ _0564_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6707 VPWR comp0.B\[0\] _0564_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X6708 _0215_ _0564_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X6709 _0564_/a_150_297# _0175_ _0564_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6710 acc0.A\[1\] _1047_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6711 _1047_/a_891_413# _1047_/a_193_47# _1047_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X6712 _1047_/a_561_413# _1047_/a_27_47# _1047_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X6713 VPWR net133 _1047_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X6714 acc0.A\[1\] _1047_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6715 _1047_/a_381_47# _0145_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X6716 VGND _1047_/a_634_159# _1047_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X6717 VPWR _1047_/a_891_413# _1047_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6718 _1047_/a_466_413# _1047_/a_193_47# _1047_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6719 VPWR _1047_/a_634_159# _1047_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6720 _1047_/a_634_159# _1047_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X6721 _1047_/a_634_159# _1047_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X6722 _1047_/a_975_413# _1047_/a_193_47# _1047_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X6723 VGND _1047_/a_1059_315# _1047_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X6724 _1047_/a_193_47# _1047_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X6725 _1047_/a_891_413# _1047_/a_27_47# _1047_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6726 _1047_/a_592_47# _1047_/a_193_47# _1047_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X6727 VPWR _1047_/a_1059_315# _1047_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6728 _1047_/a_1017_47# _1047_/a_27_47# _1047_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X6729 _1047_/a_193_47# _1047_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X6730 _1047_/a_466_413# _1047_/a_27_47# _1047_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X6731 VGND _1047_/a_891_413# _1047_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6732 _1047_/a_381_47# _0145_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6733 VGND net133 _1047_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6734 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6735 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6736 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X6737 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X6738 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6739 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6740 net121 clknet_1_1__leaf__0463_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X6741 VGND clknet_1_1__leaf__0463_ net121 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6742 net121 clknet_1_1__leaf__0463_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6743 VPWR clknet_1_1__leaf__0463_ net121 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6744 net135 clknet_1_0__leaf__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X6745 VGND clknet_1_0__leaf__0464_ net135 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6746 net135 clknet_1_0__leaf__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6747 VPWR clknet_1_0__leaf__0464_ net135 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6748 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6749 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6750 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6751 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6752 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6753 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6754 _0616_/a_78_199# _0247_ _0616_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.5655 ps=5.64 w=0.65 l=0.15
X6755 VPWR _0240_ _0616_/a_493_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X6756 _0616_/a_493_297# _0246_ _0616_/a_78_199# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.47 ps=2.94 w=1 l=0.15
X6757 VPWR _0616_/a_78_199# _0248_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.28 ps=2.56 w=1 l=0.15
X6758 VGND _0246_ _0616_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6759 _0616_/a_78_199# _0241_ _0616_/a_292_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.235 ps=2.47 w=1 l=0.15
X6760 _0616_/a_215_47# _0240_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6761 _0616_/a_215_47# _0241_ _0616_/a_78_199# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6762 _0616_/a_292_297# _0247_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6763 VGND _0616_/a_78_199# _0248_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6764 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6765 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6766 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6767 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6768 VGND comp0.B\[8\] _0547_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6769 _0547_/a_68_297# _0176_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6770 _0206_ _0547_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6771 VPWR comp0.B\[8\] _0547_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X6772 _0206_ _0547_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X6773 _0547_/a_150_297# _0176_ _0547_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6774 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6775 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6776 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6777 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6778 net116 clknet_1_1__leaf__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X6779 VGND clknet_1_1__leaf__0462_ net116 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6780 net116 clknet_1_1__leaf__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6781 VPWR clknet_1_1__leaf__0462_ net116 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6782 VPWR _0950_/a_75_212# _0161_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X6783 _0950_/a_75_212# _0469_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X6784 _0950_/a_75_212# _0469_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X6785 VGND _0950_/a_75_212# _0161_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X6786 VPWR clknet_0__0459_ clkbuf_1_1__f__0459_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X6787 VPWR clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X6788 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6789 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6790 VPWR clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6791 VPWR clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6792 clkbuf_1_1__f__0459_/a_110_47# clknet_0__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6793 clkbuf_1_1__f__0459_/a_110_47# clknet_0__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X6794 VGND clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X6795 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6796 VGND clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6797 clkbuf_1_1__f__0459_/a_110_47# clknet_0__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6798 VGND clknet_0__0459_ clkbuf_1_1__f__0459_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6799 VGND clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6800 VPWR clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6801 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6802 VGND clknet_0__0459_ clkbuf_1_1__f__0459_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6803 VGND clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6804 VPWR clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6805 VGND clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6806 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6807 clkbuf_1_1__f__0459_/a_110_47# clknet_0__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6808 VPWR clknet_0__0459_ clkbuf_1_1__f__0459_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6809 VPWR clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6810 VPWR clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6811 VGND clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6812 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6813 VGND clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6814 VGND clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6815 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6816 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6817 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6818 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6819 VPWR clkbuf_1_1__f__0459_/a_110_47# clknet_1_1__leaf__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6820 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6821 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6822 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6823 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6824 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6825 clknet_1_1__leaf__0459_ clkbuf_1_1__f__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6826 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X6827 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X6828 VPWR input19/a_75_212# net19 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X6829 input19/a_75_212# B[11] VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X6830 input19/a_75_212# B[11] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X6831 VGND input19/a_75_212# net19 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X6832 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6833 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6834 _0795_/a_81_21# _0346_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X6835 _0795_/a_299_297# _0346_ _0795_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X6836 VPWR _0795_/a_81_21# _0410_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X6837 VPWR _0405_ _0795_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6838 VGND _0795_/a_81_21# _0410_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6839 VGND _0409_ _0795_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X6840 _0795_/a_299_297# _0409_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6841 _0795_/a_384_47# _0405_ _0795_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6842 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X6843 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X6844 VPWR _0183_ _0580_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X6845 _0580_/a_27_297# _0217_ _0580_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X6846 VGND _0183_ _0580_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X6847 _0117_ _0580_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6848 _0580_/a_27_297# _0217_ _0580_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X6849 _0580_/a_109_297# acc0.A\[19\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6850 _0580_/a_373_47# acc0.A\[19\] _0580_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6851 _0117_ _0580_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6852 _0580_/a_109_297# net206 _0580_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6853 _0580_/a_109_47# net206 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6854 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6855 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6856 control0.state\[1\] _1063_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6857 _1063_/a_891_413# _1063_/a_193_47# _1063_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X6858 _1063_/a_561_413# _1063_/a_27_47# _1063_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X6859 VPWR clknet_1_1__leaf_clk _1063_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X6860 control0.state\[1\] _1063_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6861 _1063_/a_381_47# _0161_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X6862 VGND _1063_/a_634_159# _1063_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X6863 VPWR _1063_/a_891_413# _1063_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6864 _1063_/a_466_413# _1063_/a_193_47# _1063_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6865 VPWR _1063_/a_634_159# _1063_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6866 _1063_/a_634_159# _1063_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X6867 _1063_/a_634_159# _1063_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X6868 _1063_/a_975_413# _1063_/a_193_47# _1063_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X6869 VGND _1063_/a_1059_315# _1063_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X6870 _1063_/a_193_47# _1063_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X6871 _1063_/a_891_413# _1063_/a_27_47# _1063_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6872 _1063_/a_592_47# _1063_/a_193_47# _1063_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X6873 VPWR _1063_/a_1059_315# _1063_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6874 _1063_/a_1017_47# _1063_/a_27_47# _1063_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X6875 _1063_/a_193_47# _1063_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X6876 _1063_/a_466_413# _1063_/a_27_47# _1063_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X6877 VGND _1063_/a_891_413# _1063_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6878 _1063_/a_381_47# _0161_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6879 VGND clknet_1_1__leaf_clk _1063_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6880 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6881 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6882 VGND _0218_ _0778_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X6883 _0778_/a_68_297# net44 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6884 _0396_ _0778_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6885 VPWR _0218_ _0778_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X6886 _0396_ _0778_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X6887 _0778_/a_150_297# net44 _0778_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6888 VPWR _0263_ _0847_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X6889 VGND _0263_ _0450_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6890 _0847_/a_109_297# _0267_ _0450_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X6891 _0450_ _0267_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6892 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X6893 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X6894 VPWR acc0.A\[26\] hold8/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6895 VGND hold8/a_285_47# hold8/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X6896 net155 hold8/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6897 VGND acc0.A\[26\] hold8/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6898 VPWR hold8/a_285_47# hold8/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X6899 hold8/a_285_47# hold8/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X6900 hold8/a_285_47# hold8/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X6901 net155 hold8/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6902 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X6903 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X6904 VPWR _0701_/a_80_21# _0333_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X6905 _0701_/a_209_297# _0330_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.65 pd=5.3 as=0 ps=0 w=1 l=0.15
X6906 _0701_/a_303_47# _0329_ _0701_/a_209_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.208 ps=1.94 w=0.65 l=0.15
X6907 _0701_/a_209_47# _0330_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6908 VGND _0701_/a_80_21# _0333_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.17225 ps=1.83 w=0.65 l=0.15
X6909 VGND _0332_ _0701_/a_80_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2145 ps=1.96 w=0.65 l=0.15
X6910 _0701_/a_80_21# _0327_ _0701_/a_303_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6911 VPWR _0329_ _0701_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6912 _0701_/a_80_21# _0332_ _0701_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0 ps=0 w=1 l=0.15
X6913 _0701_/a_209_297# _0327_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6914 _0563_/a_240_47# net24 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X6915 _0131_ _0563_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X6916 VGND _0208_ _0563_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6917 _0563_/a_51_297# net203 _0563_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X6918 _0563_/a_149_47# _0214_ _0563_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X6919 _0563_/a_240_47# _0173_ _0563_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6920 VPWR _0208_ _0563_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X6921 _0131_ _0563_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X6922 _0563_/a_149_47# net203 _0563_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6923 _0563_/a_245_297# _0173_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6924 VPWR _0214_ _0563_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6925 _0563_/a_512_297# net24 _0563_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6926 VPWR net149 _0264_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6927 _0264_ net149 _0632_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X6928 _0632_/a_113_47# net36 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6929 _0264_ net36 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6930 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X6931 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X6932 VPWR _0494_/a_27_47# _0174_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6933 _0174_ _0494_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6934 VPWR _0173_ _0494_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X6935 _0174_ _0494_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X6936 VGND _0494_/a_27_47# _0174_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6937 VGND _0173_ _0494_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6938 comp0.B\[14\] _1046_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6939 _1046_/a_891_413# _1046_/a_193_47# _1046_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X6940 _1046_/a_561_413# _1046_/a_27_47# _1046_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X6941 VPWR net132 _1046_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X6942 comp0.B\[14\] _1046_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6943 _1046_/a_381_47# net158 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X6944 VGND _1046_/a_634_159# _1046_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X6945 VPWR _1046_/a_891_413# _1046_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6946 _1046_/a_466_413# _1046_/a_193_47# _1046_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6947 VPWR _1046_/a_634_159# _1046_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6948 _1046_/a_634_159# _1046_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X6949 _1046_/a_634_159# _1046_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X6950 _1046_/a_975_413# _1046_/a_193_47# _1046_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X6951 VGND _1046_/a_1059_315# _1046_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X6952 _1046_/a_193_47# _1046_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X6953 _1046_/a_891_413# _1046_/a_27_47# _1046_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6954 _1046_/a_592_47# _1046_/a_193_47# _1046_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X6955 VPWR _1046_/a_1059_315# _1046_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6956 _1046_/a_1017_47# _1046_/a_27_47# _1046_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X6957 _1046_/a_193_47# _1046_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X6958 _1046_/a_466_413# _1046_/a_27_47# _1046_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X6959 VGND _1046_/a_891_413# _1046_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X6960 _1046_/a_381_47# net158 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6961 VGND net132 _1046_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X6962 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X6963 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X6964 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X6965 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X6966 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X6967 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X6968 _0546_/a_240_47# net32 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X6969 _0139_ _0546_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X6970 VGND _0172_ _0546_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6971 _0546_/a_51_297# net152 _0546_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X6972 _0546_/a_149_47# _0205_ _0546_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X6973 _0546_/a_240_47# _0174_ _0546_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6974 VPWR _0172_ _0546_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X6975 _0139_ _0546_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X6976 _0546_/a_149_47# net152 _0546_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6977 _0546_/a_245_297# _0174_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6978 VPWR _0205_ _0546_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6979 _0546_/a_512_297# net32 _0546_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X6980 VPWR _0242_ _0615_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X6981 VGND _0242_ _0247_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X6982 _0615_/a_109_297# _0244_ _0247_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X6983 _0247_ _0244_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X6984 acc0.A\[29\] _1029_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X6985 _1029_/a_891_413# _1029_/a_193_47# _1029_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X6986 _1029_/a_561_413# _1029_/a_27_47# _1029_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X6987 VPWR net115 _1029_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X6988 acc0.A\[29\] _1029_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X6989 _1029_/a_381_47# net191 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X6990 VGND _1029_/a_634_159# _1029_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X6991 VPWR _1029_/a_891_413# _1029_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X6992 _1029_/a_466_413# _1029_/a_193_47# _1029_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6993 VPWR _1029_/a_634_159# _1029_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X6994 _1029_/a_634_159# _1029_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X6995 _1029_/a_634_159# _1029_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X6996 _1029_/a_975_413# _1029_/a_193_47# _1029_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X6997 VGND _1029_/a_1059_315# _1029_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X6998 _1029_/a_193_47# _1029_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X6999 _1029_/a_891_413# _1029_/a_27_47# _1029_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7000 _1029_/a_592_47# _1029_/a_193_47# _1029_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7001 VPWR _1029_/a_1059_315# _1029_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7002 _1029_/a_1017_47# _1029_/a_27_47# _1029_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7003 _1029_/a_193_47# _1029_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7004 _1029_/a_466_413# _1029_/a_27_47# _1029_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7005 VGND _1029_/a_891_413# _1029_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7006 _1029_/a_381_47# net191 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7007 VGND net115 _1029_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7008 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7009 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7010 VPWR net10 _0529_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X7011 _0529_/a_27_297# _0186_ _0529_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X7012 VGND net10 _0529_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X7013 _0197_ _0529_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7014 _0529_/a_27_297# _0186_ _0529_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X7015 _0529_/a_109_297# _0180_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7016 _0529_/a_373_47# _0180_ _0529_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7017 _0197_ _0529_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7018 _0529_/a_109_297# net170 _0529_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7019 _0529_/a_109_47# net170 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7020 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7021 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7022 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7023 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7024 VPWR clknet_1_0__leaf__0457_ _0880_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X7025 _0460_ _0880_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X7026 _0460_ _0880_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X7027 VGND clknet_1_0__leaf__0457_ _0880_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X7028 VPWR clknet_0__0458_ clkbuf_1_1__f__0458_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X7029 VPWR clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X7030 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7031 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7032 VPWR clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7033 VPWR clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7034 clkbuf_1_1__f__0458_/a_110_47# clknet_0__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7035 clkbuf_1_1__f__0458_/a_110_47# clknet_0__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X7036 VGND clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X7037 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7038 VGND clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7039 clkbuf_1_1__f__0458_/a_110_47# clknet_0__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7040 VGND clknet_0__0458_ clkbuf_1_1__f__0458_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7041 VGND clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7042 VPWR clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7043 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7044 VGND clknet_0__0458_ clkbuf_1_1__f__0458_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7045 VGND clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7046 VPWR clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7047 VGND clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7048 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7049 clkbuf_1_1__f__0458_/a_110_47# clknet_0__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7050 VPWR clknet_0__0458_ clkbuf_1_1__f__0458_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7051 VPWR clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7052 VPWR clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7053 VGND clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7054 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7055 VGND clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7056 VGND clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7057 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7058 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7059 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7060 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7061 VPWR clkbuf_1_1__f__0458_/a_110_47# clknet_1_1__leaf__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7062 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7063 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7064 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7065 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7066 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7067 clknet_1_1__leaf__0458_ clkbuf_1_1__f__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7068 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7069 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7070 net94 clknet_1_1__leaf__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7071 VGND clknet_1_1__leaf__0460_ net94 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7072 net94 clknet_1_1__leaf__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7073 VPWR clknet_1_1__leaf__0460_ net94 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7074 _0794_/a_110_297# _0297_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.265 ps=2.53 w=1 l=0.15
X7075 VGND _0297_ _0794_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.17225 ps=1.83 w=0.65 l=0.15
X7076 _0409_ _0404_ _0794_/a_110_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.105 ps=1.21 w=1 l=0.15
X7077 VPWR _0300_ _0409_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X7078 _0794_/a_27_47# _0404_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X7079 _0794_/a_326_47# _0300_ _0794_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.12675 ps=1.04 w=0.65 l=0.15
X7080 _0409_ _0277_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.635 pd=3.27 as=0.195 ps=1.39 w=1 l=0.15
X7081 _0409_ _0277_ _0794_/a_326_47# VGND sky130_fd_pr__nfet_01v8 ad=0.39325 pd=2.51 as=0.06825 ps=0.86 w=0.65 l=0.15
X7082 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7083 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7084 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7085 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7086 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7087 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7088 control0.state\[0\] _1062_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7089 _1062_/a_891_413# _1062_/a_193_47# _1062_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7090 _1062_/a_561_413# _1062_/a_27_47# _1062_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7091 VPWR clknet_1_1__leaf_clk _1062_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7092 control0.state\[0\] _1062_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7093 _1062_/a_381_47# _0160_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7094 VGND _1062_/a_634_159# _1062_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7095 VPWR _1062_/a_891_413# _1062_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7096 _1062_/a_466_413# _1062_/a_193_47# _1062_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7097 VPWR _1062_/a_634_159# _1062_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7098 _1062_/a_634_159# _1062_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7099 _1062_/a_634_159# _1062_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7100 _1062_/a_975_413# _1062_/a_193_47# _1062_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7101 VGND _1062_/a_1059_315# _1062_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7102 _1062_/a_193_47# _1062_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7103 _1062_/a_891_413# _1062_/a_27_47# _1062_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7104 _1062_/a_592_47# _1062_/a_193_47# _1062_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7105 VPWR _1062_/a_1059_315# _1062_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7106 _1062_/a_1017_47# _1062_/a_27_47# _1062_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7107 _1062_/a_193_47# _1062_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7108 _1062_/a_466_413# _1062_/a_27_47# _1062_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7109 VGND _1062_/a_891_413# _1062_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7110 _1062_/a_381_47# _0160_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7111 VGND clknet_1_1__leaf_clk _1062_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7112 _0846_/a_240_47# net233 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X7113 _0083_ _0846_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X7114 VGND _0219_ _0846_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7115 _0846_/a_51_297# _0449_ _0846_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X7116 _0846_/a_149_47# _0345_ _0846_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X7117 _0846_/a_240_47# _0448_ _0846_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7118 VPWR _0219_ _0846_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X7119 _0083_ _0846_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X7120 _0846_/a_149_47# _0449_ _0846_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7121 _0846_/a_245_297# _0448_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7122 VPWR _0345_ _0846_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7123 _0846_/a_512_297# net233 _0846_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7124 _0777_/a_377_297# _0309_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=2.42 as=0 ps=0 w=1 l=0.15
X7125 _0777_/a_47_47# _0394_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7126 _0777_/a_129_47# _0394_ _0777_/a_47_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.72 as=0.169 ps=1.82 w=0.65 l=0.15
X7127 _0777_/a_285_47# _0394_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X7128 _0395_ _0777_/a_47_47# _0777_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X7129 VGND _0309_ _0777_/a_129_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7130 VPWR _0309_ _0777_/a_47_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7131 VPWR _0777_/a_47_47# _0395_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.33 ps=2.66 w=1 l=0.15
X7132 _0395_ _0394_ _0777_/a_377_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7133 _0777_/a_285_47# _0309_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7134 VPWR _0125_ hold9/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7135 VGND hold9/a_285_47# hold9/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X7136 net156 hold9/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7137 VGND _0125_ hold9/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7138 VPWR hold9/a_285_47# hold9/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X7139 hold9/a_285_47# hold9/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X7140 hold9/a_285_47# hold9/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X7141 net156 hold9/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7142 VPWR _0221_ _0332_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7143 _0332_ _0221_ _0700_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X7144 _0700_/a_113_47# _0331_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7145 _0332_ _0331_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7146 VPWR _0261_ _0631_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X7147 VGND _0261_ _0263_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7148 _0631_/a_109_297# _0262_ _0263_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X7149 _0263_ _0262_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7150 VGND net201 _0562_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X7151 _0562_/a_68_297# _0175_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7152 _0214_ _0562_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7153 VPWR net201 _0562_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X7154 _0214_ _0562_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X7155 _0562_/a_150_297# _0175_ _0562_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7156 VPWR _0171_ _0173_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7157 _0173_ _0171_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7158 VPWR control0.sh _0173_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7159 _0493_/a_27_47# control0.sh VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7160 _0493_/a_27_47# _0171_ _0173_ VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7161 _0173_ _0171_ _0493_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7162 _0173_ control0.sh VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7163 VGND control0.sh _0493_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7164 comp0.B\[13\] _1045_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7165 _1045_/a_891_413# _1045_/a_193_47# _1045_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7166 _1045_/a_561_413# _1045_/a_27_47# _1045_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7167 VPWR net131 _1045_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7168 comp0.B\[13\] _1045_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7169 _1045_/a_381_47# net184 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7170 VGND _1045_/a_634_159# _1045_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7171 VPWR _1045_/a_891_413# _1045_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7172 _1045_/a_466_413# _1045_/a_193_47# _1045_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7173 VPWR _1045_/a_634_159# _1045_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7174 _1045_/a_634_159# _1045_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7175 _1045_/a_634_159# _1045_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7176 _1045_/a_975_413# _1045_/a_193_47# _1045_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7177 VGND _1045_/a_1059_315# _1045_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7178 _1045_/a_193_47# _1045_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7179 _1045_/a_891_413# _1045_/a_27_47# _1045_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7180 _1045_/a_592_47# _1045_/a_193_47# _1045_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7181 VPWR _1045_/a_1059_315# _1045_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7182 _1045_/a_1017_47# _1045_/a_27_47# _1045_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7183 _1045_/a_193_47# _1045_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7184 _1045_/a_466_413# _1045_/a_27_47# _1045_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7185 VGND _1045_/a_891_413# _1045_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7186 _1045_/a_381_47# net184 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7187 VGND net131 _1045_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7188 _0437_ _0435_ _0829_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.348 pd=2.78 as=0.21 ps=2.42 w=1 l=0.15
X7189 VPWR _0436_ _0437_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.7 l=0.15
X7190 _0829_/a_27_47# _0435_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X7191 _0437_ _0436_ _0829_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7192 _0829_/a_109_297# _0429_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7193 VGND _0429_ _0829_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7194 _0246_ _0614_/a_29_53# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X7195 _0614_/a_111_297# _0245_ _0614_/a_29_53# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.26 as=0.1092 ps=1.36 w=0.42 l=0.15
X7196 _0246_ _0614_/a_29_53# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X7197 _0614_/a_183_297# _0244_ _0614_/a_111_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1386 pd=1.5 as=0 ps=0 w=0.42 l=0.15
X7198 VPWR _0243_ _0614_/a_183_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7199 _0614_/a_29_53# _0244_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2226 pd=2.74 as=0 ps=0 w=0.42 l=0.15
X7200 VGND _0245_ _0614_/a_29_53# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7201 VGND _0243_ _0614_/a_29_53# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7202 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7203 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7204 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7205 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7206 VGND comp0.B\[9\] _0545_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X7207 _0545_/a_68_297# _0176_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7208 _0205_ _0545_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7209 VPWR comp0.B\[9\] _0545_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X7210 _0205_ _0545_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X7211 _0545_/a_150_297# _0176_ _0545_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7212 acc0.A\[28\] _1028_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7213 _1028_/a_891_413# _1028_/a_193_47# _1028_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7214 _1028_/a_561_413# _1028_/a_27_47# _1028_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7215 VPWR net114 _1028_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7216 acc0.A\[28\] _1028_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7217 _1028_/a_381_47# _0126_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7218 VGND _1028_/a_634_159# _1028_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7219 VPWR _1028_/a_891_413# _1028_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7220 _1028_/a_466_413# _1028_/a_193_47# _1028_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7221 VPWR _1028_/a_634_159# _1028_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7222 _1028_/a_634_159# _1028_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7223 _1028_/a_634_159# _1028_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7224 _1028_/a_975_413# _1028_/a_193_47# _1028_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7225 VGND _1028_/a_1059_315# _1028_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7226 _1028_/a_193_47# _1028_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7227 _1028_/a_891_413# _1028_/a_27_47# _1028_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7228 _1028_/a_592_47# _1028_/a_193_47# _1028_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7229 VPWR _1028_/a_1059_315# _1028_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7230 _1028_/a_1017_47# _1028_/a_27_47# _1028_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7231 _1028_/a_193_47# _1028_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7232 _1028_/a_466_413# _1028_/a_27_47# _1028_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7233 VGND _1028_/a_891_413# _1028_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7234 _1028_/a_381_47# _0126_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7235 VGND net114 _1028_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7236 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7237 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7238 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7239 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7240 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X7241 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X7242 _0528_/a_81_21# _0196_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X7243 _0528_/a_299_297# _0196_ _0528_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X7244 VPWR _0528_/a_81_21# _0148_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X7245 VPWR net170 _0528_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7246 VGND _0528_/a_81_21# _0148_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7247 VGND _0195_ _0528_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X7248 _0528_/a_299_297# _0195_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7249 _0528_/a_384_47# net170 _0528_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7250 VPWR clknet_0__0457_ clkbuf_1_1__f__0457_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X7251 VPWR clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X7252 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7253 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7254 VPWR clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7255 VPWR clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7256 clkbuf_1_1__f__0457_/a_110_47# clknet_0__0457_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7257 clkbuf_1_1__f__0457_/a_110_47# clknet_0__0457_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X7258 VGND clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X7259 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7260 VGND clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7261 clkbuf_1_1__f__0457_/a_110_47# clknet_0__0457_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7262 VGND clknet_0__0457_ clkbuf_1_1__f__0457_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7263 VGND clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7264 VPWR clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7265 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7266 VGND clknet_0__0457_ clkbuf_1_1__f__0457_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7267 VGND clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7268 VPWR clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7269 VGND clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7270 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7271 clkbuf_1_1__f__0457_/a_110_47# clknet_0__0457_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7272 VPWR clknet_0__0457_ clkbuf_1_1__f__0457_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7273 VPWR clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7274 VPWR clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7275 VGND clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7276 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7277 VGND clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7278 VGND clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7279 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7280 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7281 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7282 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7283 VPWR clkbuf_1_1__f__0457_/a_110_47# clknet_1_1__leaf__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7284 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7285 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7286 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7287 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7288 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7289 clknet_1_1__leaf__0457_ clkbuf_1_1__f__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7290 net107 clknet_1_0__leaf__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7291 VGND clknet_1_0__leaf__0461_ net107 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7292 net107 clknet_1_0__leaf__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7293 VPWR clknet_1_0__leaf__0461_ net107 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7294 _0793_/a_240_47# net42 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X7295 _0095_ _0793_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X7296 VGND _0219_ _0793_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7297 _0793_/a_51_297# _0408_ _0793_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X7298 _0793_/a_149_47# _0345_ _0793_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X7299 _0793_/a_240_47# _0407_ _0793_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7300 VPWR _0219_ _0793_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X7301 _0095_ _0793_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X7302 _0793_/a_149_47# _0408_ _0793_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7303 _0793_/a_245_297# _0407_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7304 VPWR _0345_ _0793_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7305 _0793_/a_512_297# net42 _0793_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7306 VPWR _0459_ clkbuf_0__0459_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X7307 VPWR clkbuf_0__0459_/a_110_47# clknet_0__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X7308 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7309 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7310 VPWR clkbuf_0__0459_/a_110_47# clknet_0__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7311 VPWR clkbuf_0__0459_/a_110_47# clknet_0__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7312 clkbuf_0__0459_/a_110_47# _0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7313 clkbuf_0__0459_/a_110_47# _0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X7314 VGND clkbuf_0__0459_/a_110_47# clknet_0__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X7315 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7316 VGND clkbuf_0__0459_/a_110_47# clknet_0__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7317 clkbuf_0__0459_/a_110_47# _0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7318 VGND _0459_ clkbuf_0__0459_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7319 VGND clkbuf_0__0459_/a_110_47# clknet_0__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7320 VPWR clkbuf_0__0459_/a_110_47# clknet_0__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7321 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7322 VGND _0459_ clkbuf_0__0459_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7323 VGND clkbuf_0__0459_/a_110_47# clknet_0__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7324 VPWR clkbuf_0__0459_/a_110_47# clknet_0__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7325 VGND clkbuf_0__0459_/a_110_47# clknet_0__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7326 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7327 clkbuf_0__0459_/a_110_47# _0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7328 VPWR _0459_ clkbuf_0__0459_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7329 VPWR clkbuf_0__0459_/a_110_47# clknet_0__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7330 VPWR clkbuf_0__0459_/a_110_47# clknet_0__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7331 VGND clkbuf_0__0459_/a_110_47# clknet_0__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7332 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7333 VGND clkbuf_0__0459_/a_110_47# clknet_0__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7334 VGND clkbuf_0__0459_/a_110_47# clknet_0__0459_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7335 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7336 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7337 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7338 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7339 VPWR clkbuf_0__0459_/a_110_47# clknet_0__0459_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7340 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7341 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7342 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7343 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7344 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7345 clknet_0__0459_ clkbuf_0__0459_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7346 net98 clknet_1_1__leaf__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7347 VGND clknet_1_1__leaf__0461_ net98 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7348 net98 clknet_1_1__leaf__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7349 VPWR clknet_1_1__leaf__0461_ net98 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7350 acc0.A\[15\] _1061_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7351 VPWR _1061_/a_1059_315# acc0.A\[15\] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7352 _1061_/a_891_413# _1061_/a_193_47# _1061_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X7353 _1061_/a_561_413# _1061_/a_27_47# _1061_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X7354 VPWR net147 _1061_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X7355 acc0.A\[15\] _1061_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7356 _1061_/a_381_47# _0159_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X7357 VGND _1061_/a_634_159# _1061_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7358 VGND _1061_/a_1059_315# acc0.A\[15\] VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X7359 VPWR _1061_/a_891_413# _1061_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X7360 _1061_/a_466_413# _1061_/a_193_47# _1061_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X7361 VPWR _1061_/a_634_159# _1061_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.17887 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X7362 _1061_/a_634_159# _1061_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X7363 _1061_/a_634_159# _1061_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.17887 ps=1.26 w=0.75 l=0.15
X7364 _1061_/a_975_413# _1061_/a_193_47# _1061_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X7365 VGND _1061_/a_1059_315# _1061_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X7366 _1061_/a_193_47# _1061_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X7367 _1061_/a_891_413# _1061_/a_27_47# _1061_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X7368 _1061_/a_592_47# _1061_/a_193_47# _1061_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X7369 VPWR _1061_/a_1059_315# _1061_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X7370 _1061_/a_1017_47# _1061_/a_27_47# _1061_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X7371 _1061_/a_193_47# _1061_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X7372 _1061_/a_466_413# _1061_/a_27_47# _1061_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X7373 VGND _1061_/a_891_413# _1061_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7374 _1061_/a_381_47# _0159_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X7375 VGND net147 _1061_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7376 _0449_ _0350_ _0845_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.19825 ps=1.26 w=0.65 l=0.15
X7377 _0449_ _0447_ _0845_/a_193_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3925 pd=1.785 as=0.135 ps=1.27 w=1 l=0.15
X7378 _0845_/a_193_297# _0446_ _0845_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7379 VGND _0446_ _0845_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7380 VPWR _0350_ _0449_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.3925 ps=1.785 w=1 l=0.15
X7381 _0845_/a_109_47# _0447_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.19825 pd=1.26 as=0.08775 ps=0.92 w=0.65 l=0.15
X7382 _0845_/a_109_297# _0261_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7383 _0845_/a_109_47# _0261_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X7384 _0394_ _0308_ _0776_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.348 pd=2.78 as=0.21 ps=2.42 w=1 l=0.15
X7385 VPWR _0306_ _0394_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.7 l=0.15
X7386 _0776_/a_27_47# _0308_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X7387 _0394_ _0306_ _0776_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7388 _0776_/a_109_297# _0387_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7389 VGND _0387_ _0776_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7390 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7391 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7392 net132 clknet_1_1__leaf__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7393 VGND clknet_1_1__leaf__0464_ net132 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7394 net132 clknet_1_1__leaf__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7395 VPWR clknet_1_1__leaf__0464_ net132 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7396 net146 clknet_1_1__leaf__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7397 VGND clknet_1_1__leaf__0465_ net146 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7398 net146 clknet_1_1__leaf__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7399 VPWR clknet_1_1__leaf__0465_ net146 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7400 _0561_/a_240_47# net25 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X7401 _0132_ _0561_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X7402 VGND _0208_ _0561_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7403 _0561_/a_51_297# net185 _0561_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X7404 _0561_/a_149_47# _0213_ _0561_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X7405 _0561_/a_240_47# _0173_ _0561_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7406 VPWR _0208_ _0561_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X7407 _0132_ _0561_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X7408 _0561_/a_149_47# net185 _0561_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7409 _0561_/a_245_297# _0173_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7410 VPWR _0213_ _0561_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7411 _0561_/a_512_297# net25 _0561_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7412 VPWR _0492_/a_27_47# _0172_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7413 _0172_ _0492_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7414 VPWR _0171_ _0492_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7415 _0172_ _0492_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X7416 VGND _0492_/a_27_47# _0172_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7417 VGND _0171_ _0492_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7418 VPWR acc0.A\[2\] _0630_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X7419 VGND acc0.A\[2\] _0262_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7420 _0630_/a_109_297# net58 _0262_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X7421 _0262_ net58 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7422 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X7423 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X7424 comp0.B\[12\] _1044_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7425 _1044_/a_891_413# _1044_/a_193_47# _1044_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7426 _1044_/a_561_413# _1044_/a_27_47# _1044_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7427 VPWR net130 _1044_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7428 comp0.B\[12\] _1044_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7429 _1044_/a_381_47# net194 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7430 VGND _1044_/a_634_159# _1044_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7431 VPWR _1044_/a_891_413# _1044_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7432 _1044_/a_466_413# _1044_/a_193_47# _1044_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7433 VPWR _1044_/a_634_159# _1044_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7434 _1044_/a_634_159# _1044_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7435 _1044_/a_634_159# _1044_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7436 _1044_/a_975_413# _1044_/a_193_47# _1044_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7437 VGND _1044_/a_1059_315# _1044_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7438 _1044_/a_193_47# _1044_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7439 _1044_/a_891_413# _1044_/a_27_47# _1044_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7440 _1044_/a_592_47# _1044_/a_193_47# _1044_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7441 VPWR _1044_/a_1059_315# _1044_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7442 _1044_/a_1017_47# _1044_/a_27_47# _1044_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7443 _1044_/a_193_47# _1044_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7444 _1044_/a_466_413# _1044_/a_27_47# _1044_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7445 VGND _1044_/a_891_413# _1044_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7446 _1044_/a_381_47# net194 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7447 VGND net130 _1044_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7448 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X7449 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X7450 net79 clknet_1_1__leaf__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7451 VGND clknet_1_1__leaf__0459_ net79 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7452 net79 clknet_1_1__leaf__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7453 VPWR clknet_1_1__leaf__0459_ net79 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7454 VPWR _0226_ _0381_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7455 _0381_ _0226_ _0759_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X7456 _0759_/a_113_47# _0373_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7457 _0381_ _0373_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7458 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7459 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7460 _0828_/a_199_47# _0429_ _0436_ VGND sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.182 ps=1.86 w=0.65 l=0.15
X7461 _0828_/a_113_297# _0435_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.545 pd=5.09 as=0 ps=0 w=1 l=0.15
X7462 _0436_ _0343_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7463 VPWR _0429_ _0828_/a_113_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7464 _0828_/a_113_297# _0343_ _0436_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X7465 VGND _0435_ _0828_/a_199_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7466 net72 clknet_1_1__leaf__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7467 VGND clknet_1_1__leaf__0458_ net72 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7468 net72 clknet_1_1__leaf__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7469 VPWR clknet_1_1__leaf__0458_ net72 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7470 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7471 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7472 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X7473 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X7474 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7475 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7476 VPWR acc0.A\[18\] _0613_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X7477 VGND acc0.A\[18\] _0245_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7478 _0613_/a_109_297# net45 _0245_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X7479 _0245_ net45 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7480 _0544_/a_240_47# net18 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X7481 _0140_ _0544_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X7482 VGND _0172_ _0544_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7483 _0544_/a_51_297# net198 _0544_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X7484 _0544_/a_149_47# _0204_ _0544_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X7485 _0544_/a_240_47# _0174_ _0544_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7486 VPWR _0172_ _0544_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X7487 _0140_ _0544_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X7488 _0544_/a_149_47# net198 _0544_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7489 _0544_/a_245_297# _0174_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7490 VPWR _0204_ _0544_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7491 _0544_/a_512_297# net18 _0544_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7492 net113 clknet_1_1__leaf__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7493 VGND clknet_1_1__leaf__0462_ net113 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7494 net113 clknet_1_1__leaf__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7495 VPWR clknet_1_1__leaf__0462_ net113 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7496 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7497 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7498 acc0.A\[27\] _1027_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7499 _1027_/a_891_413# _1027_/a_193_47# _1027_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7500 _1027_/a_561_413# _1027_/a_27_47# _1027_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7501 VPWR net113 _1027_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7502 acc0.A\[27\] _1027_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7503 _1027_/a_381_47# net156 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7504 VGND _1027_/a_634_159# _1027_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7505 VPWR _1027_/a_891_413# _1027_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7506 _1027_/a_466_413# _1027_/a_193_47# _1027_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7507 VPWR _1027_/a_634_159# _1027_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7508 _1027_/a_634_159# _1027_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7509 _1027_/a_634_159# _1027_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7510 _1027_/a_975_413# _1027_/a_193_47# _1027_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7511 VGND _1027_/a_1059_315# _1027_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7512 _1027_/a_193_47# _1027_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7513 _1027_/a_891_413# _1027_/a_27_47# _1027_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7514 _1027_/a_592_47# _1027_/a_193_47# _1027_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7515 VPWR _1027_/a_1059_315# _1027_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7516 _1027_/a_1017_47# _1027_/a_27_47# _1027_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7517 _1027_/a_193_47# _1027_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7518 _1027_/a_466_413# _1027_/a_27_47# _1027_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7519 VGND _1027_/a_891_413# _1027_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7520 _1027_/a_381_47# net156 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7521 VGND net113 _1027_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7522 VPWR net53 hold90/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7523 VGND hold90/a_285_47# hold90/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X7524 net237 hold90/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7525 VGND net53 hold90/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7526 VPWR hold90/a_285_47# hold90/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X7527 hold90/a_285_47# hold90/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X7528 hold90/a_285_47# hold90/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X7529 net237 hold90/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7530 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X7531 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X7532 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7533 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7534 VPWR net11 _0527_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X7535 _0527_/a_27_297# _0186_ _0527_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X7536 VGND net11 _0527_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X7537 _0196_ _0527_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7538 _0527_/a_27_297# _0186_ _0527_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X7539 _0527_/a_109_297# _0180_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7540 _0527_/a_373_47# _0180_ _0527_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7541 _0196_ _0527_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7542 _0527_/a_109_297# net154 _0527_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7543 _0527_/a_109_47# net154 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7544 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7545 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7546 VPWR _0792_/a_80_21# _0408_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X7547 _0792_/a_209_297# _0405_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.65 pd=5.3 as=0 ps=0 w=1 l=0.15
X7548 _0792_/a_303_47# _0400_ _0792_/a_209_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2145 pd=1.96 as=0.208 ps=1.94 w=0.65 l=0.15
X7549 _0792_/a_209_47# _0405_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7550 VGND _0792_/a_80_21# _0408_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.17225 ps=1.83 w=0.65 l=0.15
X7551 VGND _0343_ _0792_/a_80_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2145 ps=1.96 w=0.65 l=0.15
X7552 _0792_/a_80_21# _0406_ _0792_/a_303_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7553 VPWR _0400_ _0792_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7554 _0792_/a_80_21# _0343_ _0792_/a_209_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0 ps=0 w=1 l=0.15
X7555 _0792_/a_209_297# _0406_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7556 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X7557 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X7558 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7559 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7560 VPWR _0458_ clkbuf_0__0458_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X7561 VPWR clkbuf_0__0458_/a_110_47# clknet_0__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X7562 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7563 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7564 VPWR clkbuf_0__0458_/a_110_47# clknet_0__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7565 VPWR clkbuf_0__0458_/a_110_47# clknet_0__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7566 clkbuf_0__0458_/a_110_47# _0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7567 clkbuf_0__0458_/a_110_47# _0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X7568 VGND clkbuf_0__0458_/a_110_47# clknet_0__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X7569 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7570 VGND clkbuf_0__0458_/a_110_47# clknet_0__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7571 clkbuf_0__0458_/a_110_47# _0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7572 VGND _0458_ clkbuf_0__0458_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7573 VGND clkbuf_0__0458_/a_110_47# clknet_0__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7574 VPWR clkbuf_0__0458_/a_110_47# clknet_0__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7575 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7576 VGND _0458_ clkbuf_0__0458_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7577 VGND clkbuf_0__0458_/a_110_47# clknet_0__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7578 VPWR clkbuf_0__0458_/a_110_47# clknet_0__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7579 VGND clkbuf_0__0458_/a_110_47# clknet_0__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7580 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7581 clkbuf_0__0458_/a_110_47# _0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7582 VPWR _0458_ clkbuf_0__0458_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7583 VPWR clkbuf_0__0458_/a_110_47# clknet_0__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7584 VPWR clkbuf_0__0458_/a_110_47# clknet_0__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7585 VGND clkbuf_0__0458_/a_110_47# clknet_0__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7586 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7587 VGND clkbuf_0__0458_/a_110_47# clknet_0__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7588 VGND clkbuf_0__0458_/a_110_47# clknet_0__0458_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7589 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7590 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7591 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7592 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7593 VPWR clkbuf_0__0458_/a_110_47# clknet_0__0458_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7594 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7595 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7596 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7597 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7598 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7599 clknet_0__0458_ clkbuf_0__0458_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7600 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7601 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7602 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7603 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7604 acc0.A\[14\] _1060_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7605 _1060_/a_891_413# _1060_/a_193_47# _1060_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7606 _1060_/a_561_413# _1060_/a_27_47# _1060_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7607 VPWR net146 _1060_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7608 acc0.A\[14\] _1060_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7609 _1060_/a_381_47# _0158_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7610 VGND _1060_/a_634_159# _1060_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7611 VPWR _1060_/a_891_413# _1060_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7612 _1060_/a_466_413# _1060_/a_193_47# _1060_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7613 VPWR _1060_/a_634_159# _1060_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7614 _1060_/a_634_159# _1060_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7615 _1060_/a_634_159# _1060_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7616 _1060_/a_975_413# _1060_/a_193_47# _1060_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7617 VGND _1060_/a_1059_315# _1060_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7618 _1060_/a_193_47# _1060_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7619 _1060_/a_891_413# _1060_/a_27_47# _1060_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7620 _1060_/a_592_47# _1060_/a_193_47# _1060_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7621 VPWR _1060_/a_1059_315# _1060_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7622 _1060_/a_1017_47# _1060_/a_27_47# _1060_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7623 _1060_/a_193_47# _1060_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7624 _1060_/a_466_413# _1060_/a_27_47# _1060_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7625 VGND _1060_/a_891_413# _1060_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7626 _1060_/a_381_47# _0158_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7627 VGND net146 _1060_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7628 VPWR _0261_ _0844_/a_382_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.305 ps=2.61 w=1 l=0.15
X7629 _0844_/a_297_47# _0447_ _0844_/a_79_21# VGND sky130_fd_pr__nfet_01v8 ad=0.3705 pd=3.74 as=0.169 ps=1.82 w=0.65 l=0.15
X7630 _0844_/a_297_47# _0261_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7631 VGND _0446_ _0844_/a_297_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7632 VPWR _0844_/a_79_21# _0448_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.28 ps=2.56 w=1 l=0.15
X7633 _0844_/a_79_21# _0447_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.15
X7634 _0844_/a_382_297# _0446_ _0844_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7635 VGND _0844_/a_79_21# _0448_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7636 VPWR clknet_1_1__leaf__0457_ _0913_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.2054 ps=2.1 w=0.79 l=0.15
X7637 _0463_ _0913_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0 ps=0 w=0.52 l=0.15
X7638 _0463_ _0913_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0 ps=0 w=0.79 l=0.15
X7639 VGND clknet_1_1__leaf__0457_ _0913_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1352 ps=1.56 w=0.52 l=0.15
X7640 VGND _0347_ _0775_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X7641 _0775_/a_510_47# _0393_ _0775_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X7642 _0775_/a_79_21# _0352_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X7643 VPWR _0393_ _0775_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7644 _0775_/a_79_21# _0392_ _0775_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X7645 _0775_/a_297_297# _0347_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7646 _0775_/a_79_21# _0352_ _0775_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X7647 VPWR _0775_/a_79_21# _0098_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X7648 VGND _0775_/a_79_21# _0098_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7649 _0775_/a_215_47# _0392_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7650 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7651 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7652 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X7653 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X7654 _0171_ control0.reset VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7655 VGND control0.reset _0171_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7656 _0171_ control0.reset VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7657 VPWR control0.reset _0171_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7658 VGND comp0.B\[2\] _0560_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X7659 _0560_/a_68_297# _0175_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7660 _0213_ _0560_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7661 VPWR comp0.B\[2\] _0560_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X7662 _0213_ _0560_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X7663 _0560_/a_150_297# _0175_ _0560_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7664 comp0.B\[11\] _1043_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7665 _1043_/a_891_413# _1043_/a_193_47# _1043_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7666 _1043_/a_561_413# _1043_/a_27_47# _1043_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7667 VPWR net129 _1043_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7668 comp0.B\[11\] _1043_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7669 _1043_/a_381_47# net196 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7670 VGND _1043_/a_634_159# _1043_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7671 VPWR _1043_/a_891_413# _1043_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7672 _1043_/a_466_413# _1043_/a_193_47# _1043_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7673 VPWR _1043_/a_634_159# _1043_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7674 _1043_/a_634_159# _1043_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7675 _1043_/a_634_159# _1043_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7676 _1043_/a_975_413# _1043_/a_193_47# _1043_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7677 VGND _1043_/a_1059_315# _1043_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7678 _1043_/a_193_47# _1043_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7679 _1043_/a_891_413# _1043_/a_27_47# _1043_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7680 _1043_/a_592_47# _1043_/a_193_47# _1043_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7681 VPWR _1043_/a_1059_315# _1043_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7682 _1043_/a_1017_47# _1043_/a_27_47# _1043_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7683 _1043_/a_193_47# _1043_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7684 _1043_/a_466_413# _1043_/a_27_47# _1043_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7685 VGND _1043_/a_891_413# _1043_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7686 _1043_/a_381_47# net196 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7687 VGND net129 _1043_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7688 _0435_ _0434_ _0827_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.348 pd=2.78 as=0.21 ps=2.42 w=1 l=0.15
X7689 VPWR _0273_ _0435_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.7 l=0.15
X7690 _0827_/a_27_47# _0434_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X7691 _0435_ _0273_ _0827_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7692 _0827_/a_109_297# _0430_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7693 VGND _0430_ _0827_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7694 VGND _0347_ _0758_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X7695 _0758_/a_510_47# _0380_ _0758_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X7696 _0758_/a_79_21# _0352_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X7697 VPWR _0380_ _0758_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7698 _0758_/a_79_21# _0379_ _0758_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X7699 _0758_/a_297_297# _0347_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7700 _0758_/a_79_21# _0352_ _0758_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X7701 VPWR _0758_/a_79_21# _0102_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X7702 VGND _0758_/a_79_21# _0102_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7703 _0758_/a_215_47# _0379_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7704 VGND _0319_ _0689_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X7705 _0689_/a_68_297# _0320_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7706 _0321_ _0689_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7707 VPWR _0319_ _0689_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X7708 _0321_ _0689_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X7709 _0689_/a_150_297# _0320_ _0689_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7710 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7711 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7712 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X7713 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X7714 VPWR net45 _0612_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X7715 _0244_ _0612_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X7716 VGND net45 _0612_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X7717 _0612_/a_59_75# acc0.A\[18\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7718 _0244_ _0612_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X7719 _0612_/a_145_75# acc0.A\[18\] _0612_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X7720 VGND net152 _0543_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X7721 _0543_/a_68_297# _0176_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7722 _0204_ _0543_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7723 VPWR net152 _0543_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X7724 _0204_ _0543_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X7725 _0543_/a_150_297# _0176_ _0543_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7726 acc0.A\[26\] _1026_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7727 _1026_/a_891_413# _1026_/a_193_47# _1026_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7728 _1026_/a_561_413# _1026_/a_27_47# _1026_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7729 VPWR net112 _1026_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7730 acc0.A\[26\] _1026_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7731 _1026_/a_381_47# _0124_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7732 VGND _1026_/a_634_159# _1026_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7733 VPWR _1026_/a_891_413# _1026_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7734 _1026_/a_466_413# _1026_/a_193_47# _1026_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7735 VPWR _1026_/a_634_159# _1026_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7736 _1026_/a_634_159# _1026_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7737 _1026_/a_634_159# _1026_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7738 _1026_/a_975_413# _1026_/a_193_47# _1026_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7739 VGND _1026_/a_1059_315# _1026_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7740 _1026_/a_193_47# _1026_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7741 _1026_/a_891_413# _1026_/a_27_47# _1026_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7742 _1026_/a_592_47# _1026_/a_193_47# _1026_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7743 VPWR _1026_/a_1059_315# _1026_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7744 _1026_/a_1017_47# _1026_/a_27_47# _1026_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7745 _1026_/a_193_47# _1026_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7746 _1026_/a_466_413# _1026_/a_27_47# _1026_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7747 VGND _1026_/a_891_413# _1026_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7748 _1026_/a_381_47# _0124_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7749 VGND net112 _1026_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7750 VPWR net57 hold80/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7751 VGND hold80/a_285_47# hold80/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X7752 net227 hold80/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7753 VGND net57 hold80/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7754 VPWR hold80/a_285_47# hold80/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X7755 hold80/a_285_47# hold80/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X7756 hold80/a_285_47# hold80/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X7757 net227 hold80/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7758 VPWR net41 hold91/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7759 VGND hold91/a_285_47# hold91/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X7760 net238 hold91/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7761 VGND net41 hold91/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7762 VPWR hold91/a_285_47# hold91/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X7763 hold91/a_285_47# hold91/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X7764 hold91/a_285_47# hold91/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X7765 net238 hold91/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7766 VPWR _0178_ _0526_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X7767 VGND _0526_/a_27_47# _0195_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X7768 VGND _0526_/a_27_47# _0195_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7769 _0195_ _0526_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X7770 _0195_ _0526_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7771 VGND _0178_ _0526_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X7772 VPWR _0526_/a_27_47# _0195_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7773 _0195_ _0526_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7774 _0195_ _0526_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7775 VPWR _0526_/a_27_47# _0195_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7776 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7777 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7778 net55 _1009_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7779 _1009_/a_891_413# _1009_/a_193_47# _1009_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7780 _1009_/a_561_413# _1009_/a_27_47# _1009_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7781 VPWR net95 _1009_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7782 net55 _1009_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7783 _1009_/a_381_47# _0107_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7784 VGND _1009_/a_634_159# _1009_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7785 VPWR _1009_/a_891_413# _1009_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7786 _1009_/a_466_413# _1009_/a_193_47# _1009_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7787 VPWR _1009_/a_634_159# _1009_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7788 _1009_/a_634_159# _1009_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7789 _1009_/a_634_159# _1009_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7790 _1009_/a_975_413# _1009_/a_193_47# _1009_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7791 VGND _1009_/a_1059_315# _1009_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7792 _1009_/a_193_47# _1009_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7793 _1009_/a_891_413# _1009_/a_27_47# _1009_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7794 _1009_/a_592_47# _1009_/a_193_47# _1009_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7795 VPWR _1009_/a_1059_315# _1009_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7796 _1009_/a_1017_47# _1009_/a_27_47# _1009_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7797 _1009_/a_193_47# _1009_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7798 _1009_/a_466_413# _1009_/a_27_47# _1009_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7799 VGND _1009_/a_891_413# _1009_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7800 _1009_/a_381_47# _0107_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7801 VGND net95 _1009_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7802 net105 clknet_1_0__leaf__0461_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7803 VGND clknet_1_0__leaf__0461_ net105 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7804 net105 clknet_1_0__leaf__0461_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7805 VPWR clknet_1_0__leaf__0461_ net105 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7806 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7807 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7808 VPWR _0509_/a_27_47# _0186_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7809 _0186_ _0509_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7810 VPWR _0182_ _0509_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7811 _0186_ _0509_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X7812 VGND _0509_/a_27_47# _0186_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7813 VGND _0182_ _0509_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7814 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X7815 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X7816 _0791_/a_199_47# _0400_ _0407_ VGND sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.182 ps=1.86 w=0.65 l=0.15
X7817 _0791_/a_113_297# _0405_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.545 pd=5.09 as=0 ps=0 w=1 l=0.15
X7818 _0407_ _0406_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7819 VPWR _0400_ _0791_/a_113_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7820 _0791_/a_113_297# _0406_ _0407_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X7821 VGND _0405_ _0791_/a_199_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7822 net86 clknet_1_0__leaf__0459_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7823 VGND clknet_1_0__leaf__0459_ net86 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7824 net86 clknet_1_0__leaf__0459_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7825 VPWR clknet_1_0__leaf__0459_ net86 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7826 net65 _0989_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7827 _0989_/a_891_413# _0989_/a_193_47# _0989_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7828 _0989_/a_561_413# _0989_/a_27_47# _0989_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7829 VPWR net75 _0989_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7830 net65 _0989_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7831 _0989_/a_381_47# _0087_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7832 VGND _0989_/a_634_159# _0989_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7833 VPWR _0989_/a_891_413# _0989_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7834 _0989_/a_466_413# _0989_/a_193_47# _0989_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7835 VPWR _0989_/a_634_159# _0989_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7836 _0989_/a_634_159# _0989_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7837 _0989_/a_634_159# _0989_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7838 _0989_/a_975_413# _0989_/a_193_47# _0989_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7839 VGND _0989_/a_1059_315# _0989_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7840 _0989_/a_193_47# _0989_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7841 _0989_/a_891_413# _0989_/a_27_47# _0989_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7842 _0989_/a_592_47# _0989_/a_193_47# _0989_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7843 VPWR _0989_/a_1059_315# _0989_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7844 _0989_/a_1017_47# _0989_/a_27_47# _0989_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7845 _0989_/a_193_47# _0989_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7846 _0989_/a_466_413# _0989_/a_27_47# _0989_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7847 VGND _0989_/a_891_413# _0989_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7848 _0989_/a_381_47# _0087_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7849 VGND net75 _0989_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7850 VPWR _0457_ clkbuf_0__0457_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.56 ps=5.12 w=1 l=0.15
X7851 VPWR clkbuf_0__0457_/a_110_47# clknet_0__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=2.24 ps=20.48 w=1 l=0.15
X7852 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7853 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7854 VPWR clkbuf_0__0457_/a_110_47# clknet_0__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7855 VPWR clkbuf_0__0457_/a_110_47# clknet_0__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7856 clkbuf_0__0457_/a_110_47# _0457_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7857 clkbuf_0__0457_/a_110_47# _0457_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2352 pd=2.8 as=0 ps=0 w=0.42 l=0.15
X7858 VGND clkbuf_0__0457_/a_110_47# clknet_0__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.9408 ps=11.2 w=0.42 l=0.15
X7859 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7860 VGND clkbuf_0__0457_/a_110_47# clknet_0__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7861 clkbuf_0__0457_/a_110_47# _0457_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7862 VGND _0457_ clkbuf_0__0457_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7863 VGND clkbuf_0__0457_/a_110_47# clknet_0__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7864 VPWR clkbuf_0__0457_/a_110_47# clknet_0__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7865 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7866 VGND _0457_ clkbuf_0__0457_/a_110_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7867 VGND clkbuf_0__0457_/a_110_47# clknet_0__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7868 VPWR clkbuf_0__0457_/a_110_47# clknet_0__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7869 VGND clkbuf_0__0457_/a_110_47# clknet_0__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7870 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7871 clkbuf_0__0457_/a_110_47# _0457_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7872 VPWR _0457_ clkbuf_0__0457_/a_110_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7873 VPWR clkbuf_0__0457_/a_110_47# clknet_0__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7874 VPWR clkbuf_0__0457_/a_110_47# clknet_0__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7875 VGND clkbuf_0__0457_/a_110_47# clknet_0__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7876 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7877 VGND clkbuf_0__0457_/a_110_47# clknet_0__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7878 VGND clkbuf_0__0457_/a_110_47# clknet_0__0457_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7879 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7880 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7881 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7882 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7883 VPWR clkbuf_0__0457_/a_110_47# clknet_0__0457_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7884 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7885 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7886 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7887 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7888 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7889 clknet_0__0457_ clkbuf_0__0457_/a_110_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7890 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7891 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7892 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7893 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7894 VGND _0260_ _0843_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X7895 _0843_/a_68_297# _0268_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7896 _0447_ _0843_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7897 VPWR _0260_ _0843_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X7898 _0447_ _0843_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X7899 _0843_/a_150_297# _0268_ _0843_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7900 VGND _0218_ _0774_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X7901 _0774_/a_68_297# net45 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7902 _0393_ _0774_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7903 VPWR _0218_ _0774_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X7904 _0393_ _0774_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X7905 _0774_/a_150_297# net45 _0774_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7906 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7907 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7908 comp0.B\[10\] _1042_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7909 _1042_/a_891_413# _1042_/a_193_47# _1042_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7910 _1042_/a_561_413# _1042_/a_27_47# _1042_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7911 VPWR net128 _1042_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7912 comp0.B\[10\] _1042_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7913 _1042_/a_381_47# _0140_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7914 VGND _1042_/a_634_159# _1042_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7915 VPWR _1042_/a_891_413# _1042_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7916 _1042_/a_466_413# _1042_/a_193_47# _1042_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7917 VPWR _1042_/a_634_159# _1042_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7918 _1042_/a_634_159# _1042_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7919 _1042_/a_634_159# _1042_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7920 _1042_/a_975_413# _1042_/a_193_47# _1042_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7921 VGND _1042_/a_1059_315# _1042_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7922 _1042_/a_193_47# _1042_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7923 _1042_/a_891_413# _1042_/a_27_47# _1042_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7924 _1042_/a_592_47# _1042_/a_193_47# _1042_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7925 VPWR _1042_/a_1059_315# _1042_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7926 _1042_/a_1017_47# _1042_/a_27_47# _1042_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X7927 _1042_/a_193_47# _1042_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X7928 _1042_/a_466_413# _1042_/a_27_47# _1042_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X7929 VGND _1042_/a_891_413# _1042_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X7930 _1042_/a_381_47# _0140_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7931 VGND net128 _1042_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7932 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X7933 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X7934 _0826_/a_219_297# _0826_/a_27_53# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1575 ps=1.17 w=0.42 l=0.15
X7935 VGND _0433_ _0826_/a_27_53# VGND sky130_fd_pr__nfet_01v8 ad=0.1575 pd=1.17 as=0.1092 ps=1.36 w=0.42 l=0.15
X7936 VPWR _0255_ _0826_/a_301_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X7937 _0434_ _0826_/a_219_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.10187 ps=0.99 w=0.65 l=0.15
X7938 _0826_/a_301_297# _0826_/a_27_53# _0826_/a_219_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X7939 _0434_ _0826_/a_219_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X7940 _0826_/a_27_53# _0433_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.1092 ps=1.36 w=0.42 l=0.15
X7941 VGND _0255_ _0826_/a_219_297# VGND sky130_fd_pr__nfet_01v8 ad=0.10187 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X7942 VGND _0350_ _0757_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X7943 _0757_/a_68_297# net243 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7944 _0380_ _0757_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7945 VPWR _0350_ _0757_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X7946 _0380_ _0757_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X7947 _0757_/a_150_297# net243 _0757_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7948 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7949 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7950 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X7951 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X7952 VPWR acc0.A\[26\] _0688_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X7953 VGND acc0.A\[26\] _0320_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7954 _0688_/a_109_297# net54 _0320_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X7955 _0320_ net54 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7956 net137 clknet_1_1__leaf__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X7957 VGND clknet_1_1__leaf__0464_ net137 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X7958 net137 clknet_1_1__leaf__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7959 VPWR clknet_1_1__leaf__0464_ net137 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7960 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7961 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7962 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X7963 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X7964 _0542_/a_240_47# net19 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X7965 _0141_ _0542_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X7966 VGND _0172_ _0542_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7967 _0542_/a_51_297# net195 _0542_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X7968 _0542_/a_149_47# _0203_ _0542_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X7969 _0542_/a_240_47# _0174_ _0542_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7970 VPWR _0172_ _0542_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X7971 _0141_ _0542_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X7972 _0542_/a_149_47# net195 _0542_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X7973 _0542_/a_245_297# _0174_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7974 VPWR _0203_ _0542_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7975 _0542_/a_512_297# net19 _0542_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X7976 VGND _0241_ _0611_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X7977 _0611_/a_68_297# _0242_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7978 _0243_ _0611_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7979 VPWR _0241_ _0611_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X7980 _0243_ _0611_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X7981 _0611_/a_150_297# _0242_ _0611_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X7982 acc0.A\[25\] _1025_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X7983 _1025_/a_891_413# _1025_/a_193_47# _1025_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X7984 _1025_/a_561_413# _1025_/a_27_47# _1025_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X7985 VPWR net111 _1025_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X7986 acc0.A\[25\] _1025_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X7987 _1025_/a_381_47# net200 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X7988 VGND _1025_/a_634_159# _1025_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X7989 VPWR _1025_/a_891_413# _1025_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X7990 _1025_/a_466_413# _1025_/a_193_47# _1025_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7991 VPWR _1025_/a_634_159# _1025_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7992 _1025_/a_634_159# _1025_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X7993 _1025_/a_634_159# _1025_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X7994 _1025_/a_975_413# _1025_/a_193_47# _1025_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X7995 VGND _1025_/a_1059_315# _1025_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X7996 _1025_/a_193_47# _1025_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X7997 _1025_/a_891_413# _1025_/a_27_47# _1025_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X7998 _1025_/a_592_47# _1025_/a_193_47# _1025_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X7999 VPWR _1025_/a_1059_315# _1025_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8000 _1025_/a_1017_47# _1025_/a_27_47# _1025_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8001 _1025_/a_193_47# _1025_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8002 _1025_/a_466_413# _1025_/a_27_47# _1025_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8003 VGND _1025_/a_891_413# _1025_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8004 _1025_/a_381_47# net200 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8005 VGND net111 _1025_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8006 _0809_/a_81_21# _0289_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X8007 _0809_/a_299_297# _0289_ _0809_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X8008 VPWR _0809_/a_81_21# _0420_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X8009 VPWR _0295_ _0809_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8010 VGND _0809_/a_81_21# _0420_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8011 VGND _0401_ _0809_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X8012 _0809_/a_299_297# _0401_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8013 _0809_/a_384_47# _0295_ _0809_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8014 VPWR net37 hold70/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8015 VGND hold70/a_285_47# hold70/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8016 net217 hold70/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8017 VGND net37 hold70/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8018 VPWR hold70/a_285_47# hold70/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8019 hold70/a_285_47# hold70/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8020 hold70/a_285_47# hold70/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8021 net217 hold70/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8022 VPWR acc0.A\[12\] hold81/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8023 VGND hold81/a_285_47# hold81/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8024 net228 hold81/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8025 VGND acc0.A\[12\] hold81/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8026 VPWR hold81/a_285_47# hold81/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8027 hold81/a_285_47# hold81/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8028 hold81/a_285_47# hold81/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8029 net228 hold81/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8030 VPWR net59 hold92/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8031 VGND hold92/a_285_47# hold92/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8032 net239 hold92/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8033 VGND net59 hold92/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8034 VPWR hold92/a_285_47# hold92/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8035 hold92/a_285_47# hold92/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8036 hold92/a_285_47# hold92/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8037 net239 hold92/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8038 _0525_/a_81_21# _0194_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X8039 _0525_/a_299_297# _0194_ _0525_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X8040 VPWR _0525_/a_81_21# _0149_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X8041 VPWR net154 _0525_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8042 VGND _0525_/a_81_21# _0149_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8043 VGND _0179_ _0525_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X8044 _0525_/a_299_297# _0179_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8045 _0525_/a_384_47# net154 _0525_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8046 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8047 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8048 net54 _1008_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8049 _1008_/a_891_413# _1008_/a_193_47# _1008_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8050 _1008_/a_561_413# _1008_/a_27_47# _1008_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8051 VPWR net94 _1008_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8052 net54 _1008_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8053 _1008_/a_381_47# _0106_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8054 VGND _1008_/a_634_159# _1008_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8055 VPWR _1008_/a_891_413# _1008_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8056 _1008_/a_466_413# _1008_/a_193_47# _1008_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8057 VPWR _1008_/a_634_159# _1008_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8058 _1008_/a_634_159# _1008_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8059 _1008_/a_634_159# _1008_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8060 _1008_/a_975_413# _1008_/a_193_47# _1008_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8061 VGND _1008_/a_1059_315# _1008_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8062 _1008_/a_193_47# _1008_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8063 _1008_/a_891_413# _1008_/a_27_47# _1008_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8064 _1008_/a_592_47# _1008_/a_193_47# _1008_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8065 VPWR _1008_/a_1059_315# _1008_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8066 _1008_/a_1017_47# _1008_/a_27_47# _1008_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8067 _1008_/a_193_47# _1008_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8068 _1008_/a_466_413# _1008_/a_27_47# _1008_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8069 VGND _1008_/a_891_413# _1008_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8070 _1008_/a_381_47# _0106_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8071 VGND net94 _1008_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8072 VPWR output60/a_27_47# pp[31] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8073 pp[31] output60/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8074 VPWR net60 output60/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8075 pp[31] output60/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X8076 VGND output60/a_27_47# pp[31] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8077 VGND net60 output60/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8078 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8079 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8080 _0508_/a_81_21# _0185_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X8081 _0508_/a_299_297# _0185_ _0508_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X8082 VPWR _0508_/a_81_21# _0157_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X8083 VPWR net228 _0508_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8084 VGND _0508_/a_81_21# _0157_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8085 VGND _0179_ _0508_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X8086 _0508_/a_299_297# _0179_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8087 _0508_/a_384_47# net228 _0508_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8088 _0406_ _0790_/a_35_297# _0790_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.53 ps=5.06 w=1 l=0.15
X8089 _0406_ net42 _0790_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.5005 pd=2.84 as=0.1755 ps=1.84 w=0.65 l=0.15
X8090 _0790_/a_35_297# net42 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X8091 _0790_/a_117_297# net42 _0790_/a_35_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.26 ps=2.52 w=1 l=0.15
X8092 VPWR net42 _0790_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8093 VGND acc0.A\[15\] _0790_/a_35_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8094 VGND _0790_/a_35_297# _0406_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8095 _0790_/a_285_297# acc0.A\[15\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8096 VPWR acc0.A\[15\] _0790_/a_117_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8097 _0790_/a_285_47# acc0.A\[15\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8098 net64 _0988_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8099 _0988_/a_891_413# _0988_/a_193_47# _0988_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8100 _0988_/a_561_413# _0988_/a_27_47# _0988_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8101 VPWR net74 _0988_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8102 net64 _0988_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8103 _0988_/a_381_47# _0086_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8104 VGND _0988_/a_634_159# _0988_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8105 VPWR _0988_/a_891_413# _0988_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8106 _0988_/a_466_413# _0988_/a_193_47# _0988_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8107 VPWR _0988_/a_634_159# _0988_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8108 _0988_/a_634_159# _0988_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8109 _0988_/a_634_159# _0988_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8110 _0988_/a_975_413# _0988_/a_193_47# _0988_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8111 VGND _0988_/a_1059_315# _0988_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8112 _0988_/a_193_47# _0988_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8113 _0988_/a_891_413# _0988_/a_27_47# _0988_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8114 _0988_/a_592_47# _0988_/a_193_47# _0988_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8115 VPWR _0988_/a_1059_315# _0988_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8116 _0988_/a_1017_47# _0988_/a_27_47# _0988_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8117 _0988_/a_193_47# _0988_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8118 _0988_/a_466_413# _0988_/a_27_47# _0988_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8119 VGND _0988_/a_891_413# _0988_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8120 _0988_/a_381_47# _0086_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8121 VGND net74 _0988_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8122 net90 clknet_1_0__leaf__0460_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X8123 VGND clknet_1_0__leaf__0460_ net90 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X8124 net90 clknet_1_0__leaf__0460_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8125 VPWR clknet_1_0__leaf__0460_ net90 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8126 VPWR _0267_ _0842_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8127 _0446_ _0842_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X8128 VGND _0267_ _0842_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8129 _0842_/a_59_75# _0263_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8130 _0446_ _0842_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X8131 _0842_/a_145_75# _0263_ _0842_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X8132 _0392_ _0773_/a_35_297# _0773_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.53 ps=5.06 w=1 l=0.15
X8133 _0392_ _0388_ _0773_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.5005 pd=2.84 as=0.1755 ps=1.84 w=0.65 l=0.15
X8134 _0773_/a_35_297# _0388_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X8135 _0773_/a_117_297# _0388_ _0773_/a_35_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.26 ps=2.52 w=1 l=0.15
X8136 VPWR _0388_ _0773_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8137 VGND _0386_ _0773_/a_35_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8138 VGND _0773_/a_35_297# _0392_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8139 _0773_/a_285_297# _0386_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8140 VPWR _0386_ _0773_/a_117_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8141 _0773_/a_285_47# _0386_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8142 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8143 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8144 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8145 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8146 comp0.B\[9\] _1041_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8147 _1041_/a_891_413# _1041_/a_193_47# _1041_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8148 _1041_/a_561_413# _1041_/a_27_47# _1041_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8149 VPWR net127 _1041_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8150 comp0.B\[9\] _1041_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8151 _1041_/a_381_47# net153 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8152 VGND _1041_/a_634_159# _1041_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8153 VPWR _1041_/a_891_413# _1041_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8154 _1041_/a_466_413# _1041_/a_193_47# _1041_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8155 VPWR _1041_/a_634_159# _1041_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8156 _1041_/a_634_159# _1041_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8157 _1041_/a_634_159# _1041_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8158 _1041_/a_975_413# _1041_/a_193_47# _1041_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8159 VGND _1041_/a_1059_315# _1041_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8160 _1041_/a_193_47# _1041_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8161 _1041_/a_891_413# _1041_/a_27_47# _1041_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8162 _1041_/a_592_47# _1041_/a_193_47# _1041_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8163 VPWR _1041_/a_1059_315# _1041_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8164 _1041_/a_1017_47# _1041_/a_27_47# _1041_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8165 _1041_/a_193_47# _1041_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8166 _1041_/a_466_413# _1041_/a_27_47# _1041_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8167 VGND _1041_/a_891_413# _1041_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8168 _1041_/a_381_47# net153 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8169 VGND net127 _1041_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8170 VGND _0258_ _0825_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8171 _0825_/a_68_297# _0432_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8172 _0433_ _0825_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8173 VPWR _0258_ _0825_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X8174 _0433_ _0825_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X8175 _0825_/a_150_297# _0432_ _0825_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8176 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8177 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8178 VPWR net54 _0687_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8179 _0319_ _0687_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X8180 VGND net54 _0687_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8181 _0687_/a_59_75# acc0.A\[26\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8182 _0319_ _0687_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X8183 _0687_/a_145_75# acc0.A\[26\] _0687_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X8184 _0756_/a_377_297# _0225_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.21 pd=2.42 as=0 ps=0 w=1 l=0.15
X8185 _0756_/a_47_47# _0378_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X8186 _0756_/a_129_47# _0378_ _0756_/a_47_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.72 as=0.169 ps=1.82 w=0.65 l=0.15
X8187 _0756_/a_285_47# _0378_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.3445 pd=3.66 as=0 ps=0 w=0.65 l=0.15
X8188 _0379_ _0756_/a_47_47# _0756_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X8189 VGND _0225_ _0756_/a_129_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8190 VPWR _0225_ _0756_/a_47_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8191 VPWR _0756_/a_47_47# _0379_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.33 ps=2.66 w=1 l=0.15
X8192 _0379_ _0378_ _0756_/a_377_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8193 _0756_/a_285_47# _0225_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8194 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8195 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8196 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X8197 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X8198 VPWR net46 _0610_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8199 _0242_ _0610_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X8200 VGND net46 _0610_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8201 _0610_/a_59_75# acc0.A\[19\] VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8202 _0242_ _0610_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X8203 _0610_/a_145_75# acc0.A\[19\] _0610_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X8204 VGND comp0.B\[11\] _0541_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8205 _0541_/a_68_297# _0176_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8206 _0203_ _0541_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8207 VPWR comp0.B\[11\] _0541_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X8208 _0203_ _0541_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X8209 _0541_/a_150_297# _0176_ _0541_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8210 acc0.A\[24\] _1024_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8211 _1024_/a_891_413# _1024_/a_193_47# _1024_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8212 _1024_/a_561_413# _1024_/a_27_47# _1024_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8213 VPWR net110 _1024_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8214 acc0.A\[24\] _1024_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8215 _1024_/a_381_47# _0122_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8216 VGND _1024_/a_634_159# _1024_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8217 VPWR _1024_/a_891_413# _1024_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8218 _1024_/a_466_413# _1024_/a_193_47# _1024_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8219 VPWR _1024_/a_634_159# _1024_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8220 _1024_/a_634_159# _1024_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8221 _1024_/a_634_159# _1024_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8222 _1024_/a_975_413# _1024_/a_193_47# _1024_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8223 VGND _1024_/a_1059_315# _1024_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8224 _1024_/a_193_47# _1024_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8225 _1024_/a_891_413# _1024_/a_27_47# _1024_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8226 _1024_/a_592_47# _1024_/a_193_47# _1024_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8227 VPWR _1024_/a_1059_315# _1024_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8228 _1024_/a_1017_47# _1024_/a_27_47# _1024_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8229 _1024_/a_193_47# _1024_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8230 _1024_/a_466_413# _1024_/a_27_47# _1024_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8231 VGND _1024_/a_891_413# _1024_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8232 _1024_/a_381_47# _0122_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8233 VGND net110 _1024_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8234 _0808_/a_585_47# _0419_ _0808_/a_266_47# VGND sky130_fd_pr__nfet_01v8 ad=0.1365 pd=1.72 as=0.47125 ps=4.05 w=0.65 l=0.15
X8235 VGND _0417_ _0808_/a_266_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8236 VPWR _0808_/a_81_21# _0091_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X8237 _0808_/a_81_21# _0345_ _0808_/a_585_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8238 VGND _0808_/a_81_21# _0091_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8239 _0808_/a_266_297# _0346_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.36 pd=2.72 as=0 ps=0 w=1 l=0.15
X8240 _0808_/a_368_297# _0417_ _0808_/a_266_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.42 pd=2.84 as=0 ps=0 w=1 l=0.15
X8241 _0808_/a_266_47# _0418_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8242 _0808_/a_266_47# _0346_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8243 _0808_/a_81_21# _0418_ _0808_/a_368_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.535 pd=5.07 as=0 ps=0 w=1 l=0.15
X8244 _0808_/a_81_21# _0345_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8245 VPWR _0419_ _0808_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8246 VGND _0347_ _0739_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X8247 _0739_/a_510_47# _0365_ _0739_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X8248 _0739_/a_79_21# _0352_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X8249 VPWR _0365_ _0739_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8250 _0739_/a_79_21# _0364_ _0739_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X8251 _0739_/a_297_297# _0347_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8252 _0739_/a_79_21# _0352_ _0739_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X8253 VPWR _0739_/a_79_21# _0106_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X8254 VGND _0739_/a_79_21# _0106_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8255 _0739_/a_215_47# _0364_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8256 VPWR _0117_ hold60/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8257 VGND hold60/a_285_47# hold60/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8258 net207 hold60/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8259 VGND _0117_ hold60/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8260 VPWR hold60/a_285_47# hold60/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8261 hold60/a_285_47# hold60/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8262 hold60/a_285_47# hold60/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8263 net207 hold60/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8264 VPWR acc0.A\[1\] hold71/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8265 VGND hold71/a_285_47# hold71/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8266 net218 hold71/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8267 VGND acc0.A\[1\] hold71/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8268 VPWR hold71/a_285_47# hold71/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8269 hold71/a_285_47# hold71/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8270 hold71/a_285_47# hold71/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8271 net218 hold71/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8272 VPWR acc0.A\[13\] hold82/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8273 VGND hold82/a_285_47# hold82/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8274 net229 hold82/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8275 VGND acc0.A\[13\] hold82/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8276 VPWR hold82/a_285_47# hold82/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8277 hold82/a_285_47# hold82/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8278 hold82/a_285_47# hold82/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8279 net229 hold82/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8280 VPWR control0.state\[1\] hold93/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8281 VGND hold93/a_285_47# hold93/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8282 net240 hold93/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8283 VGND control0.state\[1\] hold93/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8284 VPWR hold93/a_285_47# hold93/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8285 hold93/a_285_47# hold93/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8286 hold93/a_285_47# hold93/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8287 net240 hold93/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8288 VPWR net12 _0524_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X8289 _0524_/a_27_297# _0186_ _0524_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X8290 VGND net12 _0524_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X8291 _0194_ _0524_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8292 _0524_/a_27_297# _0186_ _0524_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X8293 _0524_/a_109_297# _0180_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8294 _0524_/a_373_47# _0180_ _0524_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8295 _0194_ _0524_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8296 _0524_/a_109_297# net148 _0524_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8297 _0524_/a_109_47# net148 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8298 net53 _1007_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8299 _1007_/a_891_413# _1007_/a_193_47# _1007_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8300 _1007_/a_561_413# _1007_/a_27_47# _1007_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8301 VPWR net93 _1007_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8302 net53 _1007_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8303 _1007_/a_381_47# _0105_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8304 VGND _1007_/a_634_159# _1007_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8305 VPWR _1007_/a_891_413# _1007_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8306 _1007_/a_466_413# _1007_/a_193_47# _1007_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8307 VPWR _1007_/a_634_159# _1007_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8308 _1007_/a_634_159# _1007_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8309 _1007_/a_634_159# _1007_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8310 _1007_/a_975_413# _1007_/a_193_47# _1007_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8311 VGND _1007_/a_1059_315# _1007_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8312 _1007_/a_193_47# _1007_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8313 _1007_/a_891_413# _1007_/a_27_47# _1007_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8314 _1007_/a_592_47# _1007_/a_193_47# _1007_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8315 VPWR _1007_/a_1059_315# _1007_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8316 _1007_/a_1017_47# _1007_/a_27_47# _1007_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8317 _1007_/a_193_47# _1007_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8318 _1007_/a_466_413# _1007_/a_27_47# _1007_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8319 VGND _1007_/a_891_413# _1007_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8320 _1007_/a_381_47# _0105_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8321 VGND net93 _1007_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8322 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8323 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8324 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8325 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8326 VPWR output50/a_27_47# pp[22] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8327 pp[22] output50/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8328 VPWR net50 output50/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8329 pp[22] output50/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X8330 VGND output50/a_27_47# pp[22] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8331 VGND net50 output50/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8332 VPWR net61 output61/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X8333 VGND output61/a_27_47# pp[3] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X8334 VGND output61/a_27_47# pp[3] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8335 pp[3] output61/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X8336 pp[3] output61/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8337 VGND net61 output61/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X8338 VPWR output61/a_27_47# pp[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8339 pp[3] output61/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8340 pp[3] output61/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8341 VPWR output61/a_27_47# pp[3] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8342 VPWR net5 _0507_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X8343 _0507_/a_27_297# _0183_ _0507_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X8344 VGND net5 _0507_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X8345 _0185_ _0507_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8346 _0507_/a_27_297# _0183_ _0507_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X8347 _0507_/a_109_297# _0181_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8348 _0507_/a_373_47# _0181_ _0507_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8349 _0185_ _0507_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8350 _0507_/a_109_297# acc0.A\[13\] _0507_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8351 _0507_/a_109_47# acc0.A\[13\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8352 net63 _0987_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8353 _0987_/a_891_413# _0987_/a_193_47# _0987_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8354 _0987_/a_561_413# _0987_/a_27_47# _0987_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8355 VPWR net73 _0987_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8356 net63 _0987_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8357 _0987_/a_381_47# _0085_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8358 VGND _0987_/a_634_159# _0987_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8359 VPWR _0987_/a_891_413# _0987_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8360 _0987_/a_466_413# _0987_/a_193_47# _0987_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8361 VPWR _0987_/a_634_159# _0987_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8362 _0987_/a_634_159# _0987_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8363 _0987_/a_634_159# _0987_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8364 _0987_/a_975_413# _0987_/a_193_47# _0987_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8365 VGND _0987_/a_1059_315# _0987_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8366 _0987_/a_193_47# _0987_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8367 _0987_/a_891_413# _0987_/a_27_47# _0987_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8368 _0987_/a_592_47# _0987_/a_193_47# _0987_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8369 VPWR _0987_/a_1059_315# _0987_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8370 _0987_/a_1017_47# _0987_/a_27_47# _0987_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8371 _0987_/a_193_47# _0987_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8372 _0987_/a_466_413# _0987_/a_27_47# _0987_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8373 VGND _0987_/a_891_413# _0987_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8374 _0987_/a_381_47# _0085_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8375 VGND net73 _0987_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8376 net75 clknet_1_1__leaf__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X8377 VGND clknet_1_1__leaf__0458_ net75 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X8378 net75 clknet_1_1__leaf__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8379 VPWR clknet_1_1__leaf__0458_ net75 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8380 net77 clknet_1_0__leaf__0458_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X8381 VGND clknet_1_0__leaf__0458_ net77 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X8382 net77 clknet_1_0__leaf__0458_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8383 VPWR clknet_1_0__leaf__0458_ net77 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8384 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8385 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8386 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8387 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8388 VGND _0369_ _0772_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X8389 _0772_/a_510_47# _0391_ _0772_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X8390 _0772_/a_79_21# _0352_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X8391 VPWR _0391_ _0772_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8392 _0772_/a_79_21# net223 _0772_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X8393 _0772_/a_297_297# _0369_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8394 _0772_/a_79_21# _0352_ _0772_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X8395 VPWR _0772_/a_79_21# _0099_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X8396 VGND _0772_/a_79_21# _0099_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8397 _0772_/a_215_47# net223 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8398 VGND _0347_ _0841_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.455 ps=4 w=0.65 l=0.15
X8399 _0841_/a_510_47# _0445_ _0841_/a_215_47# VGND sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0 ps=0 w=0.65 l=0.15
X8400 _0841_/a_79_21# _0399_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.74 pd=5.48 as=0 ps=0 w=1 l=0.15
X8401 VPWR _0445_ _0841_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8402 _0841_/a_79_21# _0444_ _0841_/a_297_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.325 ps=2.65 w=1 l=0.15
X8403 _0841_/a_297_297# _0347_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8404 _0841_/a_79_21# _0399_ _0841_/a_510_47# VGND sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0 ps=0 w=0.65 l=0.15
X8405 VPWR _0841_/a_79_21# _0084_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X8406 VGND _0841_/a_79_21# _0084_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8407 _0841_/a_215_47# _0444_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8408 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8409 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8410 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X8411 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X8412 comp0.B\[8\] _1040_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8413 _1040_/a_891_413# _1040_/a_193_47# _1040_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8414 _1040_/a_561_413# _1040_/a_27_47# _1040_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8415 VPWR net126 _1040_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8416 comp0.B\[8\] _1040_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8417 _1040_/a_381_47# net174 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8418 VGND _1040_/a_634_159# _1040_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8419 VPWR _1040_/a_891_413# _1040_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8420 _1040_/a_466_413# _1040_/a_193_47# _1040_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8421 VPWR _1040_/a_634_159# _1040_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8422 _1040_/a_634_159# _1040_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8423 _1040_/a_634_159# _1040_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8424 _1040_/a_975_413# _1040_/a_193_47# _1040_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8425 VGND _1040_/a_1059_315# _1040_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8426 _1040_/a_193_47# _1040_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8427 _1040_/a_891_413# _1040_/a_27_47# _1040_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8428 _1040_/a_592_47# _1040_/a_193_47# _1040_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8429 VPWR _1040_/a_1059_315# _1040_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8430 _1040_/a_1017_47# _1040_/a_27_47# _1040_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8431 _1040_/a_193_47# _1040_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8432 _1040_/a_466_413# _1040_/a_27_47# _1040_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8433 VGND _1040_/a_891_413# _1040_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8434 _1040_/a_381_47# net174 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8435 VGND net126 _1040_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8436 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8437 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8438 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8439 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8440 VPWR _0271_ _0824_/a_59_75# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8441 _0432_ _0824_/a_59_75# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X8442 VGND _0271_ _0824_/a_145_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8443 _0824_/a_59_75# _0431_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8444 _0432_ _0824_/a_59_75# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X8445 _0824_/a_145_75# _0431_ _0824_/a_59_75# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1176 ps=1.4 w=0.42 l=0.15
X8446 VPWR _0227_ _0755_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X8447 VGND _0227_ _0378_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X8448 _0755_/a_109_297# _0374_ _0378_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X8449 _0378_ _0374_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8450 _0686_/a_219_297# _0686_/a_27_53# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0 ps=0 w=0.42 l=0.15
X8451 VGND _0317_ _0686_/a_27_53# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8452 VPWR _0316_ _0686_/a_301_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X8453 _0318_ _0686_/a_219_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X8454 _0686_/a_301_297# _0686_/a_27_53# _0686_/a_219_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8455 _0318_ _0686_/a_219_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X8456 _0686_/a_27_53# _0317_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0 ps=0 w=0.42 l=0.15
X8457 VGND _0316_ _0686_/a_219_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8458 net128 clknet_1_1__leaf__0464_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X8459 VGND clknet_1_1__leaf__0464_ net128 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X8460 net128 clknet_1_1__leaf__0464_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8461 VPWR clknet_1_1__leaf__0464_ net128 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8462 net142 clknet_1_1__leaf__0465_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X8463 VGND clknet_1_1__leaf__0465_ net142 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X8464 net142 clknet_1_1__leaf__0465_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8465 VPWR clknet_1_1__leaf__0465_ net142 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8466 _0540_/a_240_47# net20 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X8467 _0142_ _0540_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X8468 VGND _0172_ _0540_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8469 _0540_/a_51_297# net193 _0540_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X8470 _0540_/a_149_47# _0202_ _0540_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X8471 _0540_/a_240_47# _0174_ _0540_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8472 VPWR _0172_ _0540_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X8473 _0142_ _0540_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X8474 _0540_/a_149_47# net193 _0540_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8475 _0540_/a_245_297# _0174_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8476 VPWR _0202_ _0540_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8477 _0540_/a_512_297# net20 _0540_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8478 acc0.A\[23\] _1023_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8479 _1023_/a_891_413# _1023_/a_193_47# _1023_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8480 _1023_/a_561_413# _1023_/a_27_47# _1023_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8481 VPWR net109 _1023_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8482 acc0.A\[23\] _1023_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8483 _1023_/a_381_47# net177 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8484 VGND _1023_/a_634_159# _1023_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8485 VPWR _1023_/a_891_413# _1023_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8486 _1023_/a_466_413# _1023_/a_193_47# _1023_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8487 VPWR _1023_/a_634_159# _1023_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8488 _1023_/a_634_159# _1023_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8489 _1023_/a_634_159# _1023_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8490 _1023_/a_975_413# _1023_/a_193_47# _1023_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8491 VGND _1023_/a_1059_315# _1023_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8492 _1023_/a_193_47# _1023_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8493 _1023_/a_891_413# _1023_/a_27_47# _1023_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8494 _1023_/a_592_47# _1023_/a_193_47# _1023_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8495 VPWR _1023_/a_1059_315# _1023_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8496 _1023_/a_1017_47# _1023_/a_27_47# _1023_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8497 _1023_/a_193_47# _1023_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8498 _1023_/a_466_413# _1023_/a_27_47# _1023_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8499 VGND _1023_/a_891_413# _1023_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8500 _1023_/a_381_47# net177 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8501 VGND net109 _1023_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8502 VGND _0218_ _0807_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8503 _0807_/a_68_297# net246 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8504 _0419_ _0807_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8505 VPWR _0218_ _0807_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X8506 _0419_ _0807_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X8507 _0807_/a_150_297# net246 _0807_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8508 VGND _0350_ _0738_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8509 _0738_/a_68_297# net244 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8510 _0365_ _0738_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8511 VPWR _0350_ _0738_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X8512 _0365_ _0738_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X8513 _0738_/a_150_297# net244 _0738_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8514 _0301_ _0669_/a_29_53# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X8515 _0669_/a_111_297# _0300_ _0669_/a_29_53# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.26 as=0.1092 ps=1.36 w=0.42 l=0.15
X8516 _0301_ _0669_/a_29_53# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X8517 _0669_/a_183_297# _0277_ _0669_/a_111_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1386 pd=1.5 as=0 ps=0 w=0.42 l=0.15
X8518 VPWR _0276_ _0669_/a_183_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8519 _0669_/a_29_53# _0277_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.2226 pd=2.74 as=0 ps=0 w=0.42 l=0.15
X8520 VGND _0300_ _0669_/a_29_53# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8521 VGND _0276_ _0669_/a_29_53# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8522 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8523 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8524 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8525 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8526 VPWR acc0.A\[27\] hold50/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8527 VGND hold50/a_285_47# hold50/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8528 net197 hold50/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8529 VGND acc0.A\[27\] hold50/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8530 VPWR hold50/a_285_47# hold50/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8531 hold50/a_285_47# hold50/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8532 hold50/a_285_47# hold50/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8533 net197 hold50/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8534 VPWR acc0.A\[30\] hold61/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8535 VGND hold61/a_285_47# hold61/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8536 net208 hold61/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8537 VGND acc0.A\[30\] hold61/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8538 VPWR hold61/a_285_47# hold61/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8539 hold61/a_285_47# hold61/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8540 hold61/a_285_47# hold61/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8541 net208 hold61/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8542 VPWR acc0.A\[17\] hold72/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8543 VGND hold72/a_285_47# hold72/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8544 net219 hold72/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8545 VGND acc0.A\[17\] hold72/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8546 VPWR hold72/a_285_47# hold72/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8547 hold72/a_285_47# hold72/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8548 hold72/a_285_47# hold72/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8549 net219 hold72/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8550 VPWR acc0.A\[6\] hold83/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8551 VGND hold83/a_285_47# hold83/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8552 net230 hold83/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8553 VGND acc0.A\[6\] hold83/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8554 VPWR hold83/a_285_47# hold83/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8555 hold83/a_285_47# hold83/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8556 hold83/a_285_47# hold83/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8557 net230 hold83/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8558 VPWR net51 hold94/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8559 VGND hold94/a_285_47# hold94/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8560 net241 hold94/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8561 VGND net51 hold94/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8562 VPWR hold94/a_285_47# hold94/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8563 hold94/a_285_47# hold94/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8564 hold94/a_285_47# hold94/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8565 net241 hold94/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8566 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8567 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8568 net109 clknet_1_0__leaf__0462_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0 ps=0 w=1 l=0.15
X8569 VGND clknet_1_0__leaf__0462_ net109 VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X8570 net109 clknet_1_0__leaf__0462_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8571 VPWR clknet_1_0__leaf__0462_ net109 VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8572 _0523_/a_81_21# _0193_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X8573 _0523_/a_299_297# _0193_ _0523_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X8574 VPWR _0523_/a_81_21# _0150_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X8575 VPWR net148 _0523_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8576 VGND _0523_/a_81_21# _0150_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8577 VGND _0179_ _0523_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X8578 _0523_/a_299_297# _0179_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8579 _0523_/a_384_47# net148 _0523_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8580 net52 _1006_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8581 _1006_/a_891_413# _1006_/a_193_47# _1006_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8582 _1006_/a_561_413# _1006_/a_27_47# _1006_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8583 VPWR net92 _1006_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8584 net52 _1006_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8585 _1006_/a_381_47# _0104_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8586 VGND _1006_/a_634_159# _1006_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8587 VPWR _1006_/a_891_413# _1006_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8588 _1006_/a_466_413# _1006_/a_193_47# _1006_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8589 VPWR _1006_/a_634_159# _1006_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8590 _1006_/a_634_159# _1006_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8591 _1006_/a_634_159# _1006_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8592 _1006_/a_975_413# _1006_/a_193_47# _1006_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8593 VGND _1006_/a_1059_315# _1006_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8594 _1006_/a_193_47# _1006_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8595 _1006_/a_891_413# _1006_/a_27_47# _1006_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8596 _1006_/a_592_47# _1006_/a_193_47# _1006_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8597 VPWR _1006_/a_1059_315# _1006_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8598 _1006_/a_1017_47# _1006_/a_27_47# _1006_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8599 _1006_/a_193_47# _1006_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8600 _1006_/a_466_413# _1006_/a_27_47# _1006_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8601 VGND _1006_/a_891_413# _1006_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8602 _1006_/a_381_47# _0104_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8603 VGND net92 _1006_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8604 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8605 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8606 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X8607 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X8608 VPWR output51/a_27_47# pp[23] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8609 pp[23] output51/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8610 VPWR net51 output51/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8611 pp[23] output51/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X8612 VGND output51/a_27_47# pp[23] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8613 VGND net51 output51/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8614 VPWR output40/a_27_47# pp[13] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8615 pp[13] output40/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8616 VPWR net40 output40/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8617 pp[13] output40/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X8618 VGND output40/a_27_47# pp[13] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8619 VGND net40 output40/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8620 VPWR net62 output62/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X8621 VGND output62/a_27_47# pp[4] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X8622 VGND output62/a_27_47# pp[4] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8623 pp[4] output62/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X8624 pp[4] output62/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8625 VGND net62 output62/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X8626 VPWR output62/a_27_47# pp[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8627 pp[4] output62/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8628 pp[4] output62/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8629 VPWR output62/a_27_47# pp[4] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8630 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8631 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8632 _0506_/a_81_21# _0184_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0 ps=0 w=0.65 l=0.15
X8633 _0506_/a_299_297# _0184_ _0506_/a_81_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.54 pd=5.08 as=0.26 ps=2.52 w=1 l=0.15
X8634 VPWR _0506_/a_81_21# _0158_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X8635 VPWR net229 _0506_/a_299_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8636 VGND _0506_/a_81_21# _0158_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8637 VGND _0179_ _0506_/a_384_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.182 ps=1.86 w=0.65 l=0.15
X8638 _0506_/a_299_297# _0179_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8639 _0506_/a_384_47# net229 _0506_/a_81_21# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8640 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8641 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8642 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X8643 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X8644 net62 _0986_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8645 _0986_/a_891_413# _0986_/a_193_47# _0986_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8646 _0986_/a_561_413# _0986_/a_27_47# _0986_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8647 VPWR net72 _0986_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8648 net62 _0986_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8649 _0986_/a_381_47# _0084_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8650 VGND _0986_/a_634_159# _0986_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8651 VPWR _0986_/a_891_413# _0986_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8652 _0986_/a_466_413# _0986_/a_193_47# _0986_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8653 VPWR _0986_/a_634_159# _0986_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8654 _0986_/a_634_159# _0986_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8655 _0986_/a_634_159# _0986_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8656 _0986_/a_975_413# _0986_/a_193_47# _0986_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8657 VGND _0986_/a_1059_315# _0986_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8658 _0986_/a_193_47# _0986_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8659 _0986_/a_891_413# _0986_/a_27_47# _0986_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8660 _0986_/a_592_47# _0986_/a_193_47# _0986_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8661 VPWR _0986_/a_1059_315# _0986_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8662 _0986_/a_1017_47# _0986_/a_27_47# _0986_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8663 _0986_/a_193_47# _0986_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8664 _0986_/a_466_413# _0986_/a_27_47# _0986_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8665 VGND _0986_/a_891_413# _0986_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8666 _0986_/a_381_47# _0084_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8667 VGND net72 _0986_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8668 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8669 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8670 _0771_/a_298_297# _0771_/a_27_413# _0771_/a_215_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.535 pd=5.07 as=0.265 ps=2.53 w=1 l=0.15
X8671 _0771_/a_215_297# _0771_/a_27_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X8672 _0771_/a_298_297# _0389_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8673 _0391_ _0771_/a_215_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8674 VPWR _0390_ _0771_/a_27_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8675 _0391_ _0771_/a_215_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8676 _0771_/a_382_47# _0243_ _0771_/a_215_297# VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X8677 VGND _0390_ _0771_/a_27_413# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X8678 VPWR _0243_ _0771_/a_298_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8679 VGND _0389_ _0771_/a_382_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8680 VGND _0218_ _0840_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8681 _0840_/a_68_297# net62 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8682 _0445_ _0840_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8683 VPWR _0218_ _0840_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X8684 _0445_ _0840_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X8685 _0840_/a_150_297# net62 _0840_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8686 VPWR _0468_ _0969_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X8687 VGND _0468_ _0487_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X8688 _0969_/a_109_297# _0486_ _0487_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X8689 _0487_ _0486_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8690 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.05
X8691 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.05
X8692 _0754_/a_240_47# net241 VGND VGND sky130_fd_pr__nfet_01v8 ad=0.351 pd=3.68 as=0 ps=0 w=0.65 l=0.15
X8693 _0103_ _0754_/a_51_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0 ps=0 w=0.65 l=0.15
X8694 VGND _0219_ _0754_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8695 _0754_/a_51_297# _0377_ _0754_/a_245_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=1.165 pd=6.33 as=0.21 ps=2.42 w=1 l=0.15
X8696 _0754_/a_149_47# _0345_ _0754_/a_51_297# VGND sky130_fd_pr__nfet_01v8 ad=0.36725 pd=3.73 as=0.2015 ps=1.92 w=0.65 l=0.15
X8697 _0754_/a_240_47# _0376_ _0754_/a_149_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8698 VPWR _0219_ _0754_/a_512_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X8699 _0103_ _0754_/a_51_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0 ps=0 w=1 l=0.15
X8700 _0754_/a_149_47# _0377_ _0754_/a_240_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8701 _0754_/a_245_297# _0376_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8702 VPWR _0345_ _0754_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8703 _0754_/a_512_297# net241 _0754_/a_51_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8704 VPWR _0260_ _0823_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.21 ps=2.42 w=1 l=0.15
X8705 VGND _0260_ _0431_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1755 ps=1.84 w=0.65 l=0.15
X8706 _0823_/a_109_297# _0269_ _0431_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.26 ps=2.52 w=1 l=0.15
X8707 _0431_ _0269_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8708 VGND acc0.A\[27\] _0685_/a_68_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1134 ps=1.38 w=0.42 l=0.15
X8709 _0685_/a_68_297# net55 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8710 _0317_ _0685_/a_68_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8711 VPWR acc0.A\[27\] _0685_/a_150_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.0882 ps=1.26 w=0.42 l=0.15
X8712 _0317_ _0685_/a_68_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0 ps=0 w=1 l=0.15
X8713 _0685_/a_150_297# net55 _0685_/a_68_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8714 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X8715 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X8716 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=1.97
X8717 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=1.97
X8718 acc0.A\[22\] _1022_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8719 _1022_/a_891_413# _1022_/a_193_47# _1022_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8720 _1022_/a_561_413# _1022_/a_27_47# _1022_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8721 VPWR net108 _1022_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8722 acc0.A\[22\] _1022_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8723 _1022_/a_381_47# net151 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8724 VGND _1022_/a_634_159# _1022_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8725 VPWR _1022_/a_891_413# _1022_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8726 _1022_/a_466_413# _1022_/a_193_47# _1022_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8727 VPWR _1022_/a_634_159# _1022_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8728 _1022_/a_634_159# _1022_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8729 _1022_/a_634_159# _1022_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8730 _1022_/a_975_413# _1022_/a_193_47# _1022_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8731 VGND _1022_/a_1059_315# _1022_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8732 _1022_/a_193_47# _1022_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8733 _1022_/a_891_413# _1022_/a_27_47# _1022_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8734 _1022_/a_592_47# _1022_/a_193_47# _1022_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8735 VPWR _1022_/a_1059_315# _1022_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8736 _1022_/a_1017_47# _1022_/a_27_47# _1022_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8737 _1022_/a_193_47# _1022_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8738 _1022_/a_466_413# _1022_/a_27_47# _1022_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8739 VGND _1022_/a_891_413# _1022_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8740 _1022_/a_381_47# net151 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8741 VGND net108 _1022_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8742 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X8743 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X8744 VPWR _0297_ _0668_/a_382_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.305 ps=2.61 w=1 l=0.15
X8745 _0668_/a_297_47# _0299_ _0668_/a_79_21# VGND sky130_fd_pr__nfet_01v8 ad=0.3705 pd=3.74 as=0.169 ps=1.82 w=0.65 l=0.15
X8746 _0668_/a_297_47# _0297_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8747 VGND _0298_ _0668_/a_297_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8748 VPWR _0668_/a_79_21# _0300_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.28 ps=2.56 w=1 l=0.15
X8749 _0668_/a_79_21# _0299_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.39 pd=2.78 as=0 ps=0 w=1 l=0.15
X8750 _0668_/a_382_297# _0298_ _0668_/a_79_21# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8751 VGND _0668_/a_79_21# _0300_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8752 _0364_ _0737_/a_35_297# _0737_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.53 ps=5.06 w=1 l=0.15
X8753 _0364_ _0360_ _0737_/a_285_47# VGND sky130_fd_pr__nfet_01v8 ad=0.5005 pd=2.84 as=0.1755 ps=1.84 w=0.65 l=0.15
X8754 _0737_/a_35_297# _0360_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X8755 _0737_/a_117_297# _0360_ _0737_/a_35_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.26 ps=2.52 w=1 l=0.15
X8756 VPWR _0360_ _0737_/a_285_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8757 VGND _0321_ _0737_/a_35_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8758 VGND _0737_/a_35_297# _0364_ VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8759 _0737_/a_285_297# _0321_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8760 VPWR _0321_ _0737_/a_117_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8761 _0737_/a_285_47# _0321_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8762 _0806_/a_199_47# _0281_ _0418_ VGND sky130_fd_pr__nfet_01v8 ad=0.19175 pd=1.89 as=0.182 ps=1.86 w=0.65 l=0.15
X8763 _0806_/a_113_297# _0402_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.545 pd=5.09 as=0 ps=0 w=1 l=0.15
X8764 _0418_ _0286_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8765 VPWR _0281_ _0806_/a_113_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8766 _0806_/a_113_297# _0286_ _0418_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X8767 VGND _0402_ _0806_/a_199_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8768 VPWR acc0.A\[23\] _0231_ VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8769 _0231_ acc0.A\[23\] _0599_/a_113_47# VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1755 ps=1.84 w=0.65 l=0.15
X8770 _0599_/a_113_47# net51 VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8771 _0231_ net51 VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8772 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8773 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8774 VPWR acc0.A\[20\] hold40/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8775 VGND hold40/a_285_47# hold40/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8776 net187 hold40/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8777 VGND acc0.A\[20\] hold40/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8778 VPWR hold40/a_285_47# hold40/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8779 hold40/a_285_47# hold40/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8780 hold40/a_285_47# hold40/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8781 net187 hold40/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8782 VPWR comp0.B\[11\] hold51/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8783 VGND hold51/a_285_47# hold51/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8784 net198 hold51/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8785 VGND comp0.B\[11\] hold51/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8786 VPWR hold51/a_285_47# hold51/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8787 hold51/a_285_47# hold51/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8788 hold51/a_285_47# hold51/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8789 net198 hold51/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8790 VPWR _0128_ hold62/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8791 VGND hold62/a_285_47# hold62/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8792 net209 hold62/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8793 VGND _0128_ hold62/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8794 VPWR hold62/a_285_47# hold62/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8795 hold62/a_285_47# hold62/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8796 hold62/a_285_47# hold62/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8797 net209 hold62/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8798 VPWR net48 hold73/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8799 VGND hold73/a_285_47# hold73/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8800 net220 hold73/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8801 VGND net48 hold73/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8802 VPWR hold73/a_285_47# hold73/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8803 hold73/a_285_47# hold73/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8804 hold73/a_285_47# hold73/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8805 net220 hold73/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8806 VPWR control0.sh hold84/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8807 VGND hold84/a_285_47# hold84/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8808 net231 hold84/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8809 VGND control0.sh hold84/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8810 VPWR hold84/a_285_47# hold84/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8811 hold84/a_285_47# hold84/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8812 hold84/a_285_47# hold84/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8813 net231 hold84/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8814 VPWR net56 hold95/a_49_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8815 VGND hold95/a_285_47# hold95/a_391_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8816 net242 hold95/a_391_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8817 VGND net56 hold95/a_49_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8818 VPWR hold95/a_285_47# hold95/a_391_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.5
X8819 hold95/a_285_47# hold95/a_49_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8820 hold95/a_285_47# hold95/a_49_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.5
X8821 net242 hold95/a_391_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8822 VPWR net13 _0522_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X8823 _0522_/a_27_297# _0186_ _0522_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X8824 VGND net13 _0522_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X8825 _0193_ _0522_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8826 _0522_/a_27_297# _0186_ _0522_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X8827 _0522_/a_109_297# _0180_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8828 _0522_/a_373_47# _0180_ _0522_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8829 _0193_ _0522_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8830 _0522_/a_109_297# acc0.A\[6\] _0522_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8831 _0522_/a_109_47# acc0.A\[6\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8832 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=0.59
X8833 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=0.59
X8834 net51 _1005_/a_1059_315# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8835 _1005_/a_891_413# _1005_/a_193_47# _1005_/a_634_159# VGND sky130_fd_pr__special_nfet_01v8 ad=0.1368 pd=1.48 as=0.1978 ps=1.99 w=0.36 l=0.15
X8836 _1005_/a_561_413# _1005_/a_27_47# _1005_/a_466_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1533 pd=1.57 as=0.1365 ps=1.49 w=0.42 l=0.15
X8837 VPWR net91 _1005_/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8838 net51 _1005_/a_1059_315# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8839 _1005_/a_381_47# _0103_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=1.39 as=0 ps=0 w=0.42 l=0.15
X8840 VGND _1005_/a_634_159# _1005_/a_592_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1392 ps=1.53 w=0.42 l=0.15
X8841 VPWR _1005_/a_891_413# _1005_/a_1059_315# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8842 _1005_/a_466_413# _1005_/a_193_47# _1005_/a_381_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8843 VPWR _1005_/a_634_159# _1005_/a_561_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8844 _1005_/a_634_159# _1005_/a_466_413# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.64 l=0.15
X8845 _1005_/a_634_159# _1005_/a_466_413# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.219 pd=2.15 as=0 ps=0 w=0.75 l=0.15
X8846 _1005_/a_975_413# _1005_/a_193_47# _1005_/a_891_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1764 pd=1.68 as=0.1134 ps=1.38 w=0.42 l=0.15
X8847 VGND _1005_/a_1059_315# _1005_/a_1017_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.132 ps=1.49 w=0.42 l=0.15
X8848 _1005_/a_193_47# _1005_/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0 ps=0 w=0.42 l=0.15
X8849 _1005_/a_891_413# _1005_/a_27_47# _1005_/a_634_159# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8850 _1005_/a_592_47# _1005_/a_193_47# _1005_/a_466_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1242 ps=1.41 w=0.36 l=0.15
X8851 VPWR _1005_/a_1059_315# _1005_/a_975_413# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8852 _1005_/a_1017_47# _1005_/a_27_47# _1005_/a_891_413# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.36 l=0.15
X8853 _1005_/a_193_47# _1005_/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0 ps=0 w=0.64 l=0.15
X8854 _1005_/a_466_413# _1005_/a_27_47# _1005_/a_381_47# VGND sky130_fd_pr__special_nfet_01v8 ad=0 pd=0 as=0.1626 ps=1.66 w=0.36 l=0.15
X8855 VGND _1005_/a_891_413# _1005_/a_1059_315# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.169 ps=1.82 w=0.65 l=0.15
X8856 _1005_/a_381_47# _0103_ VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8857 VGND net91 _1005_/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8858 VPWR output52/a_27_47# pp[24] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8859 pp[24] output52/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8860 VPWR net52 output52/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8861 pp[24] output52/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X8862 VGND output52/a_27_47# pp[24] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8863 VGND net52 output52/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8864 VPWR output41/a_27_47# pp[14] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.27 ps=2.54 w=1 l=0.15
X8865 pp[14] output41/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8866 VPWR net41 output41/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.1664 ps=1.8 w=0.64 l=0.15
X8867 pp[14] output41/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0 ps=0 w=0.65 l=0.15
X8868 VGND output41/a_27_47# pp[14] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8869 VGND net41 output41/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1092 ps=1.36 w=0.42 l=0.15
X8870 VPWR net63 output63/a_27_47# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.265 ps=2.53 w=1 l=0.15
X8871 VGND output63/a_27_47# pp[5] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2352 ps=2.8 w=0.42 l=0.15
X8872 VGND output63/a_27_47# pp[5] VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8873 pp[5] output63/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.56 pd=5.12 as=0 ps=0 w=1 l=0.15
X8874 pp[5] output63/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8875 VGND net63 output63/a_27_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.1113 ps=1.37 w=0.42 l=0.15
X8876 VPWR output63/a_27_47# pp[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8877 pp[5] output63/a_27_47# VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.42 l=0.15
X8878 pp[5] output63/a_27_47# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8879 VPWR output63/a_27_47# pp[5] VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8880 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=4.73
X8881 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=4.73
X8882 VPWR VGND VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=0.87 l=2.89
X8883 VGND VPWR VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.55 l=2.89
X8884 VPWR net6 _0505_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0.59 ps=5.18 w=1 l=0.15
X8885 _0505_/a_27_297# _0183_ _0505_/a_109_47# VGND sky130_fd_pr__nfet_01v8 ad=0.338 pd=3.64 as=0.1495 ps=1.76 w=0.65 l=0.15
X8886 VGND net6 _0505_/a_373_47# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.2275 ps=2 w=0.65 l=0.15
X8887 _0184_ _0505_/a_27_297# VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0 ps=0 w=1 l=0.15
X8888 _0505_/a_27_297# _0183_ _0505_/a_109_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0.51285 pd=5.04 as=0 ps=0 w=1 l=0.15
X8889 _0505_/a_109_297# _0181_ VPWR VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8890 _0505_/a_373_47# _0181_ _0505_/a_27_297# VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
X8891 _0184_ _0505_/a_27_297# VGND VGND sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0 ps=0 w=0.65 l=0.15
X8892 _0505_/a_109_297# acc0.A\[14\] _0505_/a_27_297# VPWR sky130_fd_pr__pfet_01v8_hvt ad=0 pd=0 as=0 ps=0 w=1 l=0.15
X8893 _0505_/a_109_47# acc0.A\[14\] VGND VGND sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.65 l=0.15
