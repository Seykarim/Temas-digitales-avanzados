* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

X_15194__107 clknet_1_1__leaf__02750_ VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__inv_2
X_09671_ mapped_spi_ram.rcv_data\[27\] net17 _05362_ VGND VGND VPWR VPWR _05363_ sky130_fd_sc_hd__a21o_1
X_08622_ CPU.aluIn1\[20\] _04246_ VGND VGND VPWR VPWR _04342_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08553_ CPU.aluIn1\[7\] _04272_ VGND VGND VPWR VPWR _04273_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_124_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08484_ CPU.Bimm\[12\] net1295 VGND VGND VPWR VPWR _04204_ sky130_fd_sc_hd__and2_1
XFILLER_0_43_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09105_ _04816_ VGND VGND VPWR VPWR _04817_ sky130_fd_sc_hd__dlymetal6s2s_1
X_14653__761 clknet_1_0__leaf__02681_ VGND VGND VPWR VPWR net793 sky130_fd_sc_hd__inv_2
XFILLER_0_32_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09036_ _04734_ _04750_ VGND VGND VPWR VPWR _04751_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold340 CPU.registerFile\[5\]\[5\] VGND VGND VPWR VPWR net1581 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold351 _04145_ VGND VGND VPWR VPWR net1592 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold362 CPU.registerFile\[30\]\[21\] VGND VGND VPWR VPWR net1603 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold373 CPU.registerFile\[14\]\[22\] VGND VGND VPWR VPWR net1614 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 CPU.registerFile\[18\]\[23\] VGND VGND VPWR VPWR net1625 sky130_fd_sc_hd__dlygate4sd3_1
Xhold395 CPU.registerFile\[4\]\[7\] VGND VGND VPWR VPWR net1636 sky130_fd_sc_hd__dlygate4sd3_1
X_09938_ _05493_ net1699 _05559_ VGND VGND VPWR VPWR _05561_ sky130_fd_sc_hd__mux2_1
X_14051__327 clknet_1_0__leaf__08365_ VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__inv_2
X_09869_ _05007_ VGND VGND VPWR VPWR _05514_ sky130_fd_sc_hd__clkbuf_4
Xhold1040 CPU.registerFile\[1\]\[4\] VGND VGND VPWR VPWR net2281 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1051 CPU.registerFile\[27\]\[27\] VGND VGND VPWR VPWR net2292 sky130_fd_sc_hd__dlygate4sd3_1
X_11900_ net2148 _05679_ _06711_ VGND VGND VPWR VPWR _06716_ sky130_fd_sc_hd__mux2_1
Xhold1062 CPU.registerFile\[30\]\[7\] VGND VGND VPWR VPWR net2303 sky130_fd_sc_hd__dlygate4sd3_1
X_12880_ _07260_ VGND VGND VPWR VPWR _07322_ sky130_fd_sc_hd__buf_4
XFILLER_0_87_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1073 CPU.registerFile\[20\]\[4\] VGND VGND VPWR VPWR net2314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1084 CPU.registerFile\[21\]\[31\] VGND VGND VPWR VPWR net2325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1095 CPU.registerFile\[1\]\[26\] VGND VGND VPWR VPWR net2336 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_202 _07841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_213 _07999_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11831_ _06679_ VGND VGND VPWR VPWR _01652_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_224 clknet_1_0__leaf__02720_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_235 _02855_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_246 _03158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_257 _05050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_268 _05381_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11762_ _04731_ net2398 _06639_ VGND VGND VPWR VPWR _06643_ sky130_fd_sc_hd__mux2_1
XANTENNA_279 _05551_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13501_ CPU.registerFile\[16\]\[18\] CPU.registerFile\[20\]\[18\] _07233_ VGND VGND
+ VPWR VPWR _07926_ sky130_fd_sc_hd__mux2_1
X_10713_ _05520_ net1738 _06045_ VGND VGND VPWR VPWR _06050_ sky130_fd_sc_hd__mux2_1
X_14736__836 clknet_1_0__leaf__02689_ VGND VGND VPWR VPWR net868 sky130_fd_sc_hd__inv_2
XFILLER_0_82_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11693_ mapped_spi_ram.rcv_data\[13\] _06590_ _06599_ _06594_ VGND VGND VPWR VPWR
+ _01709_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16220_ _08397_ _03691_ _03695_ _02949_ VGND VGND VPWR VPWR _03696_ sky130_fd_sc_hd__a211o_1
X_13432_ _07330_ _07859_ VGND VGND VPWR VPWR _07860_ sky130_fd_sc_hd__or2_1
XFILLER_0_107_920 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10644_ mapped_spi_flash.rcv_data\[2\] _05969_ VGND VGND VPWR VPWR _06007_ sky130_fd_sc_hd__or2_1
X_16151_ _05010_ _03625_ _03628_ VGND VGND VPWR VPWR _03629_ sky130_fd_sc_hd__or3_2
XFILLER_0_51_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13363_ _07388_ _07792_ VGND VGND VPWR VPWR _07793_ sky130_fd_sc_hd__or2_1
X_10575_ _05966_ VGND VGND VPWR VPWR _05967_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer7 net1249 VGND VGND VPWR VPWR net1248 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_134_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15102_ per_uart.uart0.enable16_counter\[10\] _07188_ net1445 VGND VGND VPWR VPWR
+ _02738_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_122_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12314_ CPU.aluIn1\[1\] _06970_ _06859_ VGND VGND VPWR VPWR _06971_ sky130_fd_sc_hd__mux2_1
X_16082_ _02914_ _03559_ _03561_ _02864_ VGND VGND VPWR VPWR _03562_ sky130_fd_sc_hd__a211o_1
X_13294_ CPU.registerFile\[28\]\[11\] CPU.registerFile\[24\]\[11\] _07399_ VGND VGND
+ VPWR VPWR _07726_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12245_ _06918_ VGND VGND VPWR VPWR _01442_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_2_Left_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_39_Left_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12176_ CPU.aluShamt\[1\] CPU.aluShamt\[0\] VGND VGND VPWR VPWR _06866_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_75_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11127_ net2411 _05704_ _06263_ VGND VGND VPWR VPWR _06270_ sky130_fd_sc_hd__mux2_1
X_16984_ clknet_leaf_21_clk _01310_ VGND VGND VPWR VPWR CPU.rs2\[15\] sky130_fd_sc_hd__dfxtp_1
X_14782__878 clknet_1_1__leaf__02693_ VGND VGND VPWR VPWR net910 sky130_fd_sc_hd__inv_2
XFILLER_0_155_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11058_ net1712 _05704_ _06226_ VGND VGND VPWR VPWR _06233_ sky130_fd_sc_hd__mux2_1
X_15935_ _02796_ _03418_ VGND VGND VPWR VPWR _03419_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10009_ net2074 _04714_ _05596_ VGND VGND VPWR VPWR _05599_ sky130_fd_sc_hd__mux2_1
X_15866_ CPU.registerFile\[6\]\[13\] _03057_ _03140_ _03351_ VGND VGND VPWR VPWR _03352_
+ sky130_fd_sc_hd__o211a_1
X_17605_ net794 _01893_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_14817_ clknet_1_1__leaf__07222_ VGND VGND VPWR VPWR _02697_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_35_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15797_ CPU.registerFile\[6\]\[11\] _03057_ _03140_ _03284_ VGND VGND VPWR VPWR _03285_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_35_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14028__307 clknet_1_1__leaf__08362_ VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__inv_2
XFILLER_0_129_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17536_ net725 _01824_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17467_ net656 _01755_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16418_ CPU.registerFile\[31\]\[29\] _03072_ VGND VGND VPWR VPWR _03888_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17398_ net587 _01686_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16349_ CPU.registerFile\[24\]\[27\] _08403_ _02874_ _03820_ VGND VGND VPWR VPWR
+ _03821_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_95_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18019_ net1192 _02299_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15202__114 clknet_1_0__leaf__02751_ VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__inv_2
XFILLER_0_10_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09723_ _04817_ _05412_ VGND VGND VPWR VPWR _05413_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_126_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09654_ _04917_ _05346_ VGND VGND VPWR VPWR _05347_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_2_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08605_ CPU.aluIn1\[12\] _04261_ VGND VGND VPWR VPWR _04325_ sky130_fd_sc_hd__and2_1
X_09585_ _04504_ _04636_ VGND VGND VPWR VPWR _05280_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08536_ CPU.aluIn1\[15\] _04255_ VGND VGND VPWR VPWR _04256_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10360_ _05537_ net2369 _05799_ VGND VGND VPWR VPWR _05802_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09019_ _04471_ _04734_ VGND VGND VPWR VPWR _04735_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10291_ _05537_ net2516 _05762_ VGND VGND VPWR VPWR _05765_ sky130_fd_sc_hd__mux2_1
X_12030_ _04696_ net2132 _06783_ VGND VGND VPWR VPWR _06785_ sky130_fd_sc_hd__mux2_1
Xhold170 CPU.cycles\[18\] VGND VGND VPWR VPWR net1411 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold181 _07173_ VGND VGND VPWR VPWR net1422 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 CPU.cycles\[21\] VGND VGND VPWR VPWR net1433 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15720_ _03208_ _03209_ _08400_ VGND VGND VPWR VPWR _03210_ sky130_fd_sc_hd__mux2_1
X_12932_ _07262_ VGND VGND VPWR VPWR _07373_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15651_ _02821_ VGND VGND VPWR VPWR _03143_ sky130_fd_sc_hd__clkbuf_4
X_12863_ _07305_ VGND VGND VPWR VPWR _07306_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_158_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11814_ _05381_ net1956 _06661_ VGND VGND VPWR VPWR _06670_ sky130_fd_sc_hd__mux2_1
X_18370_ net38 net29 VGND VGND VPWR VPWR mapped_spi_ram.div_counter\[2\] sky130_fd_sc_hd__dfxtp_1
X_15582_ _03072_ _03073_ _03075_ VGND VGND VPWR VPWR _03076_ sky130_fd_sc_hd__o21a_1
X_12794_ _04936_ _05336_ VGND VGND VPWR VPWR _07237_ sky130_fd_sc_hd__nand2_2
XFILLER_0_157_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17321_ net510 _01609_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14324__465 clknet_1_0__leaf__08465_ VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__inv_2
XFILLER_0_68_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11745_ net1344 _06627_ _06630_ _06632_ VGND VGND VPWR VPWR _01691_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17252_ net442 _01540_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_13962__247 clknet_1_1__leaf__08356_ VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__inv_2
XFILLER_0_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11676_ _06574_ VGND VGND VPWR VPWR _06590_ sky130_fd_sc_hd__buf_2
XFILLER_0_154_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_670 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16203_ _03671_ _03678_ _05361_ VGND VGND VPWR VPWR _03679_ sky130_fd_sc_hd__mux2_1
X_13415_ CPU.registerFile\[2\]\[15\] CPU.registerFile\[3\]\[15\] _07263_ VGND VGND
+ VPWR VPWR _07843_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17183_ clknet_leaf_25_clk _01471_ VGND VGND VPWR VPWR CPU.Jimm\[13\] sky130_fd_sc_hd__dfxtp_2
X_10627_ mapped_spi_flash.rcv_data\[10\] _05994_ VGND VGND VPWR VPWR _05998_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_40_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16134_ CPU.registerFile\[27\]\[21\] CPU.registerFile\[31\]\[21\] _08403_ VGND VGND
+ VPWR VPWR _03612_ sky130_fd_sc_hd__mux2_1
X_13346_ CPU.registerFile\[13\]\[13\] _07772_ _07773_ CPU.registerFile\[9\]\[13\]
+ _07775_ VGND VGND VPWR VPWR _07776_ sky130_fd_sc_hd__o221a_1
XFILLER_0_52_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10558_ net1430 _05950_ _05952_ _05954_ VGND VGND VPWR VPWR _02202_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_47_Left_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16065_ _03252_ _03536_ _03544_ _02935_ VGND VGND VPWR VPWR _03545_ sky130_fd_sc_hd__o211a_1
X_13277_ CPU.registerFile\[6\]\[11\] CPU.registerFile\[7\]\[11\] _07371_ VGND VGND
+ VPWR VPWR _07709_ sky130_fd_sc_hd__mux2_1
X_10489_ _04512_ net1289 _04544_ VGND VGND VPWR VPWR _05898_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12228_ _06905_ VGND VGND VPWR VPWR _01446_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_90_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14034__311 clknet_1_0__leaf__08364_ VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__inv_2
X_12159_ _06852_ VGND VGND VPWR VPWR _01496_ sky130_fd_sc_hd__clkbuf_1
X_16967_ net262 _01293_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_108_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765__215 clknet_1_0__leaf__07224_ VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__inv_2
X_15918_ CPU.registerFile\[9\]\[15\] CPU.registerFile\[13\]\[15\] _02999_ VGND VGND
+ VPWR VPWR _03402_ sky130_fd_sc_hd__mux2_1
X_16898_ _06515_ VGND VGND VPWR VPWR _04176_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_56_Left_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15849_ CPU.registerFile\[8\]\[13\] _02789_ _03117_ _03334_ VGND VGND VPWR VPWR _03335_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_88_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09370_ CPU.aluIn1\[16\] _04254_ _04698_ _04808_ CPU.aluReg\[16\] VGND VGND VPWR
+ VPWR _05075_ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14719__820 clknet_1_0__leaf__02688_ VGND VGND VPWR VPWR net852 sky130_fd_sc_hd__inv_2
XFILLER_0_19_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17519_ net708 _01807_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14299__442 clknet_1_0__leaf__08463_ VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__inv_2
XFILLER_0_46_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14080__353 clknet_1_0__leaf__08368_ VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__inv_2
XFILLER_0_46_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_65_Left_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_136_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14765__862 clknet_1_0__leaf__02692_ VGND VGND VPWR VPWR net894 sky130_fd_sc_hd__inv_2
X_16525__192 clknet_1_1__leaf__03964_ VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_74_Left_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09706_ _05395_ _05396_ _04670_ VGND VGND VPWR VPWR _05397_ sky130_fd_sc_hd__mux2_1
X_09637_ _04916_ _05327_ _05329_ _04974_ _05330_ VGND VGND VPWR VPWR _05331_ sky130_fd_sc_hd__o221a_1
XFILLER_0_139_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09568_ _04671_ _05263_ VGND VGND VPWR VPWR _05264_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_26_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08519_ CPU.rs2\[22\] _04200_ _04205_ VGND VGND VPWR VPWR _04239_ sky130_fd_sc_hd__a21o_1
X_09499_ _04265_ _04740_ VGND VGND VPWR VPWR _05198_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_156_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_156_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11530_ _04589_ _06491_ VGND VGND VPWR VPWR _06492_ sky130_fd_sc_hd__nor2_2
XFILLER_0_81_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_83_Left_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_137_Right_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11461_ _06447_ VGND VGND VPWR VPWR _01793_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13200_ _07268_ _07631_ _07634_ VGND VGND VPWR VPWR _07635_ sky130_fd_sc_hd__or3_1
XFILLER_0_33_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10412_ _05830_ _05837_ VGND VGND VPWR VPWR _05838_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_59_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11392_ _05516_ net2408 _06408_ VGND VGND VPWR VPWR _06411_ sky130_fd_sc_hd__mux2_1
X_14180_ clknet_1_1__leaf__08363_ VGND VGND VPWR VPWR _08428_ sky130_fd_sc_hd__buf_1
XFILLER_0_61_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13131_ CPU.registerFile\[16\]\[7\] CPU.registerFile\[20\]\[7\] _07457_ VGND VGND
+ VPWR VPWR _07567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10343_ _05520_ net1887 _05788_ VGND VGND VPWR VPWR _05793_ sky130_fd_sc_hd__mux2_1
X_14848__937 clknet_1_0__leaf__02700_ VGND VGND VPWR VPWR net969 sky130_fd_sc_hd__inv_2
X_13062_ _07237_ VGND VGND VPWR VPWR _07500_ sky130_fd_sc_hd__clkbuf_8
X_10274_ _05520_ net2455 _05751_ VGND VGND VPWR VPWR _05756_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12013_ _06775_ VGND VGND VPWR VPWR _01566_ sky130_fd_sc_hd__clkbuf_1
X_17870_ net1059 _02154_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[28\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_92_Left_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16821_ per_uart.uart0.tx_count16\[2\] _04121_ net1593 VGND VGND VPWR VPWR _04124_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_136_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16752_ _04001_ _04067_ _04068_ _04069_ _07123_ VGND VGND VPWR VPWR _04070_ sky130_fd_sc_hd__o311a_1
XFILLER_0_45_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15703_ CPU.registerFile\[8\]\[9\] CPU.registerFile\[12\]\[9\] _02798_ VGND VGND
+ VPWR VPWR _03193_ sky130_fd_sc_hd__mux2_1
X_12915_ _07230_ _07335_ _07356_ _07309_ VGND VGND VPWR VPWR _07357_ sky130_fd_sc_hd__a211o_1
X_16683_ _08436_ _08459_ _05329_ VGND VGND VPWR VPWR _04011_ sky130_fd_sc_hd__a21o_1
X_13895_ _08305_ _08307_ _04972_ VGND VGND VPWR VPWR _08308_ sky130_fd_sc_hd__mux2_1
X_15634_ CPU.registerFile\[9\]\[7\] _02778_ _03125_ VGND VGND VPWR VPWR _03126_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12846_ _07235_ VGND VGND VPWR VPWR _07289_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_103_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14894__979 clknet_1_1__leaf__02704_ VGND VGND VPWR VPWR net1011 sky130_fd_sc_hd__inv_2
X_18353_ clknet_leaf_6_clk net1685 VGND VGND VPWR VPWR per_uart.uart0.rx_bitcount\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_15231__140 clknet_1_1__leaf__02754_ VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__inv_2
XFILLER_0_28_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15565_ CPU.registerFile\[6\]\[5\] _03057_ _02894_ _03058_ VGND VGND VPWR VPWR _03059_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17304_ net493 _01592_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18284_ net117 _02564_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_11728_ net22 _06617_ net1309 net8 VGND VGND VPWR VPWR _06620_ sky130_fd_sc_hd__a31o_1
XFILLER_0_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15496_ _02809_ _02988_ _02991_ VGND VGND VPWR VPWR _02992_ sky130_fd_sc_hd__or3_2
XFILLER_0_154_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17235_ net425 _01523_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[28\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_104_Right_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11659_ _06515_ VGND VGND VPWR VPWR _06581_ sky130_fd_sc_hd__buf_2
XFILLER_0_25_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17166_ net390 _01454_ VGND VGND VPWR VPWR CPU.aluReg\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__08431_ _08431_ VGND VGND VPWR VPWR clknet_0__08431_ sky130_fd_sc_hd__clkbuf_16
Xhold906 CPU.registerFile\[16\]\[22\] VGND VGND VPWR VPWR net2147 sky130_fd_sc_hd__dlygate4sd3_1
X_16117_ _02914_ _03593_ _03595_ _02864_ VGND VGND VPWR VPWR _03596_ sky130_fd_sc_hd__a211o_1
Xhold917 CPU.registerFile\[29\]\[4\] VGND VGND VPWR VPWR net2158 sky130_fd_sc_hd__dlygate4sd3_1
Xhold928 CPU.registerFile\[26\]\[13\] VGND VGND VPWR VPWR net2169 sky130_fd_sc_hd__dlygate4sd3_1
X_13329_ _07351_ _07759_ VGND VGND VPWR VPWR _07760_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17097_ net355 _01419_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[27\] sky130_fd_sc_hd__dfxtp_1
Xhold939 CPU.registerFile\[29\]\[3\] VGND VGND VPWR VPWR net2180 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__02755_ clknet_0__02755_ VGND VGND VPWR VPWR clknet_1_1__leaf__02755_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0__08362_ _08362_ VGND VGND VPWR VPWR clknet_0__08362_ sky130_fd_sc_hd__clkbuf_16
X_16048_ _02936_ _03521_ _03528_ _02934_ VGND VGND VPWR VPWR _03529_ sky130_fd_sc_hd__o211a_1
Xclkbuf_1_1__f__02686_ clknet_0__02686_ VGND VGND VPWR VPWR clknet_1_1__leaf__02686_
+ sky130_fd_sc_hd__clkbuf_16
X_08870_ _04589_ CPU.state\[2\] CPU.state\[3\] VGND VGND VPWR VPWR _04590_ sky130_fd_sc_hd__nor3_4
XTAP_TAPCELL_ROW_4_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17999_ clknet_leaf_7_clk _02283_ VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[13\]
+ sky130_fd_sc_hd__dfxtp_1
X_09422_ _04895_ _05124_ VGND VGND VPWR VPWR _05125_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09353_ _04442_ _04701_ VGND VGND VPWR VPWR _05059_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_23_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09284_ _04248_ _04339_ _04340_ VGND VGND VPWR VPWR _04993_ sky130_fd_sc_hd__o21a_1
XFILLER_0_90_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14006__287 clknet_1_1__leaf__08360_ VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_134_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload90 clknet_1_1__leaf__08433_ VGND VGND VPWR VPWR clkload90/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14353__491 clknet_1_1__leaf__08468_ VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_54_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__03962_ clknet_0__03962_ VGND VGND VPWR VPWR clknet_1_0__leaf__03962_
+ sky130_fd_sc_hd__clkbuf_16
X_13991__273 clknet_1_1__leaf__08359_ VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__inv_2
X_08999_ _04487_ VGND VGND VPWR VPWR _04716_ sky130_fd_sc_hd__clkbuf_4
X_10961_ net1608 _05675_ _06179_ VGND VGND VPWR VPWR _06182_ sky130_fd_sc_hd__mux2_1
X_12700_ net1339 _07181_ VGND VGND VPWR VPWR _07182_ sky130_fd_sc_hd__or2_1
X_13680_ CPU.registerFile\[4\]\[23\] _07374_ VGND VGND VPWR VPWR _08100_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10892_ _06145_ VGND VGND VPWR VPWR _02060_ sky130_fd_sc_hd__clkbuf_1
X_12631_ CPU.cycles\[4\] CPU.cycles\[5\] _07138_ VGND VGND VPWR VPWR _07140_ sky130_fd_sc_hd__and3_1
X_15350_ _05093_ VGND VGND VPWR VPWR _02848_ sky130_fd_sc_hd__buf_4
X_12562_ net2349 _05129_ _07096_ VGND VGND VPWR VPWR _07104_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11513_ net10 _06473_ VGND VGND VPWR VPWR _06478_ sky130_fd_sc_hd__and2b_1
X_15281_ _02779_ VGND VGND VPWR VPWR _02780_ sky130_fd_sc_hd__buf_4
XFILLER_0_109_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12493_ _07067_ VGND VGND VPWR VPWR _01343_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17020_ net278 _01342_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_11444_ _06438_ VGND VGND VPWR VPWR _01801_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_684 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14436__566 clknet_1_0__leaf__02659_ VGND VGND VPWR VPWR net598 sky130_fd_sc_hd__inv_2
X_14163_ _08418_ VGND VGND VPWR VPWR _01482_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11375_ _05499_ CPU.registerFile\[24\]\[27\] _06397_ VGND VGND VPWR VPWR _06402_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13114_ CPU.registerFile\[14\]\[6\] CPU.registerFile\[10\]\[6\] _07274_ VGND VGND
+ VPWR VPWR _07551_ sky130_fd_sc_hd__mux2_1
X_10326_ _05503_ CPU.registerFile\[21\]\[25\] _05777_ VGND VGND VPWR VPWR _05784_
+ sky130_fd_sc_hd__mux2_1
X_14094_ _05134_ _04621_ _08369_ VGND VGND VPWR VPWR _08374_ sky130_fd_sc_hd__o21a_1
X_13045_ CPU.registerFile\[31\]\[4\] _07482_ _07420_ CPU.registerFile\[27\]\[4\] _07483_
+ VGND VGND VPWR VPWR _07484_ sky130_fd_sc_hd__o221a_1
X_17922_ net1111 _02206_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[2\] sky130_fd_sc_hd__dfxtp_1
X_10257_ _05503_ net2377 _05740_ VGND VGND VPWR VPWR _05747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10188_ _05701_ VGND VGND VPWR VPWR _02335_ sky130_fd_sc_hd__clkbuf_1
X_17853_ net1042 _02137_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16804_ net1511 VGND VGND VPWR VPWR _04112_ sky130_fd_sc_hd__inv_2
X_17784_ net973 _02068_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_14902__986 clknet_1_0__leaf__02705_ VGND VGND VPWR VPWR net1018 sky130_fd_sc_hd__inv_2
X_16735_ _04049_ _04055_ _04015_ VGND VGND VPWR VPWR _02592_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_85_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16666_ _08457_ _03993_ _03994_ _03996_ VGND VGND VPWR VPWR _03997_ sky130_fd_sc_hd__a31o_1
X_14601__714 clknet_1_0__leaf__02676_ VGND VGND VPWR VPWR net746 sky130_fd_sc_hd__inv_2
X_13878_ CPU.registerFile\[29\]\[29\] _07289_ _07290_ CPU.registerFile\[25\]\[29\]
+ _07249_ VGND VGND VPWR VPWR _08292_ sky130_fd_sc_hd__o221a_1
XFILLER_0_76_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15617_ CPU.registerFile\[20\]\[6\] CPU.registerFile\[21\]\[6\] _02829_ VGND VGND
+ VPWR VPWR _03110_ sky130_fd_sc_hd__mux2_1
X_12829_ _05338_ VGND VGND VPWR VPWR _07272_ sky130_fd_sc_hd__buf_4
XFILLER_0_158_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_754 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15548_ CPU.registerFile\[13\]\[5\] _02775_ VGND VGND VPWR VPWR _03042_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18336_ clknet_leaf_4_clk _02616_ VGND VGND VPWR VPWR per_uart.rx_data\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18267_ clknet_leaf_1_clk _02547_ VGND VGND VPWR VPWR per_uart.uart0.rxd_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15479_ _02924_ _02972_ _02973_ _02974_ _02930_ VGND VGND VPWR VPWR _02975_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17218_ net408 _01506_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18198_ net229 _02478_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_116_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold703 CPU.registerFile\[9\]\[27\] VGND VGND VPWR VPWR net1944 sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 CPU.registerFile\[13\]\[16\] VGND VGND VPWR VPWR net1955 sky130_fd_sc_hd__dlygate4sd3_1
X_17149_ net373 _01437_ VGND VGND VPWR VPWR CPU.aluReg\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold725 CPU.registerFile\[17\]\[11\] VGND VGND VPWR VPWR net1966 sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 CPU.registerFile\[31\]\[20\] VGND VGND VPWR VPWR net1977 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold747 CPU.registerFile\[26\]\[4\] VGND VGND VPWR VPWR net1988 sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 CPU.registerFile\[23\]\[24\] VGND VGND VPWR VPWR net1999 sky130_fd_sc_hd__dlygate4sd3_1
X_09971_ _05526_ net2198 _05570_ VGND VGND VPWR VPWR _05578_ sky130_fd_sc_hd__mux2_1
Xhold769 CPU.registerFile\[17\]\[2\] VGND VGND VPWR VPWR net2010 sky130_fd_sc_hd__dlygate4sd3_1
X_08922_ _04631_ _04641_ _04635_ VGND VGND VPWR VPWR _04642_ sky130_fd_sc_hd__and3b_1
Xclkbuf_1_1__f__02669_ clknet_0__02669_ VGND VGND VPWR VPWR clknet_1_1__leaf__02669_
+ sky130_fd_sc_hd__clkbuf_16
X_08853_ CPU.aluIn1\[20\] _04495_ VGND VGND VPWR VPWR _04573_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08784_ CPU.Jimm\[13\] VGND VGND VPWR VPWR _04504_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_28_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14877__963 clknet_1_0__leaf__02703_ VGND VGND VPWR VPWR net995 sky130_fd_sc_hd__inv_2
XFILLER_0_95_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09405_ _05108_ VGND VGND VPWR VPWR _05109_ sky130_fd_sc_hd__buf_4
XFILLER_0_153_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09336_ CPU.PC\[18\] _04926_ VGND VGND VPWR VPWR _05043_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09267_ CPU.PC\[21\] _04928_ VGND VGND VPWR VPWR _04977_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09198_ CPU.PC\[22\] _04821_ _04909_ VGND VGND VPWR VPWR _04910_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11160_ _05557_ _05738_ VGND VGND VPWR VPWR _06287_ sky130_fd_sc_hd__nand2_4
XFILLER_0_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10111_ CPU.registerFile\[18\]\[13\] _05150_ _05644_ VGND VGND VPWR VPWR _05653_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11091_ _04665_ _04664_ CPU.writeBack _04663_ VGND VGND VPWR VPWR _06250_ sky130_fd_sc_hd__or4bb_4
X_10042_ net2257 _05150_ _05607_ VGND VGND VPWR VPWR _05616_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold74 _06031_ VGND VGND VPWR VPWR net1315 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 mapped_spi_ram.cmd_addr\[25\] VGND VGND VPWR VPWR net1326 sky130_fd_sc_hd__dlygate4sd3_1
X_13801_ _07650_ _08215_ _08216_ VGND VGND VPWR VPWR _08217_ sky130_fd_sc_hd__o21ai_1
Xhold96 net7 VGND VGND VPWR VPWR net1337 sky130_fd_sc_hd__dlygate4sd3_1
X_11993_ _05109_ net2405 _06758_ VGND VGND VPWR VPWR _06765_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13732_ _07268_ _08145_ _08149_ VGND VGND VPWR VPWR _08150_ sky130_fd_sc_hd__or3_1
X_10944_ _06172_ VGND VGND VPWR VPWR _02035_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_67_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16451_ CPU.registerFile\[16\]\[30\] CPU.registerFile\[18\]\[30\] _08400_ VGND VGND
+ VPWR VPWR _03920_ sky130_fd_sc_hd__mux2_1
X_13663_ CPU.registerFile\[31\]\[23\] _08082_ _07256_ CPU.registerFile\[27\]\[23\]
+ _07320_ VGND VGND VPWR VPWR _08083_ sky130_fd_sc_hd__a221o_1
X_10875_ _06135_ VGND VGND VPWR VPWR _02067_ sky130_fd_sc_hd__clkbuf_1
X_15402_ CPU.registerFile\[16\]\[1\] CPU.registerFile\[18\]\[1\] _08399_ VGND VGND
+ VPWR VPWR _02900_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__02689_ clknet_0__02689_ VGND VGND VPWR VPWR clknet_1_0__leaf__02689_
+ sky130_fd_sc_hd__clkbuf_16
X_12614_ _06479_ _07130_ VGND VGND VPWR VPWR _07131_ sky130_fd_sc_hd__or2_1
X_16382_ _02812_ _03849_ _03852_ _02948_ VGND VGND VPWR VPWR _03853_ sky130_fd_sc_hd__o211a_1
X_13594_ _06515_ VGND VGND VPWR VPWR _08017_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_80_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18121_ net184 _02401_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_14_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15333_ _02831_ VGND VGND VPWR VPWR _02832_ sky130_fd_sc_hd__clkbuf_4
X_12545_ net1679 _04957_ _07085_ VGND VGND VPWR VPWR _07095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18052_ net1225 _02332_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_15264_ _05406_ VGND VGND VPWR VPWR _02763_ sky130_fd_sc_hd__clkbuf_8
X_12476_ _07058_ VGND VGND VPWR VPWR _01351_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17003_ clknet_leaf_11_clk _00002_ VGND VGND VPWR VPWR CPU.state\[2\] sky130_fd_sc_hd__dfxtp_2
XANTENNA_5 _02787_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11427_ _05551_ CPU.registerFile\[24\]\[2\] _06419_ VGND VGND VPWR VPWR _06429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_20_Left_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14146_ _08407_ VGND VGND VPWR VPWR _08408_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11358_ _05551_ net1960 _06382_ VGND VGND VPWR VPWR _06392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10309_ _05555_ net1891 _05739_ VGND VGND VPWR VPWR _05774_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11289_ _06355_ VGND VGND VPWR VPWR _01873_ sky130_fd_sc_hd__clkbuf_1
X_17905_ net1094 _02189_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[23\] sky130_fd_sc_hd__dfxtp_2
X_13028_ _07364_ _07466_ VGND VGND VPWR VPWR _07467_ sky130_fd_sc_hd__or2_1
X_17836_ net1025 _02120_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[26\] sky130_fd_sc_hd__dfxtp_1
Xrebuffer17 net1259 VGND VGND VPWR VPWR net1258 sky130_fd_sc_hd__dlygate4sd1_1
X_17767_ net956 _02051_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[21\] sky130_fd_sc_hd__dfxtp_1
Xrebuffer28 net1270 VGND VGND VPWR VPWR net1269 sky130_fd_sc_hd__dlymetal6s2s_1
Xrebuffer39 _04532_ VGND VGND VPWR VPWR net1280 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_77_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16718_ _08379_ _05197_ _04006_ VGND VGND VPWR VPWR _04041_ sky130_fd_sc_hd__or3b_1
XFILLER_0_88_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17698_ net887 _01986_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09121_ CPU.PC\[19\] _04832_ VGND VGND VPWR VPWR _04833_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_33_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18319_ clknet_leaf_15_clk _02599_ VGND VGND VPWR VPWR CPU.PC\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09052_ _04353_ _04236_ _04351_ VGND VGND VPWR VPWR _04766_ sky130_fd_sc_hd__or3_1
XFILLER_0_32_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14419__550 clknet_1_0__leaf__02658_ VGND VGND VPWR VPWR net582 sky130_fd_sc_hd__inv_2
XFILLER_0_114_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold500 CPU.registerFile\[20\]\[18\] VGND VGND VPWR VPWR net1741 sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 CPU.registerFile\[16\]\[25\] VGND VGND VPWR VPWR net1752 sky130_fd_sc_hd__dlygate4sd3_1
Xhold522 CPU.PC\[20\] VGND VGND VPWR VPWR net1763 sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 CPU.registerFile\[17\]\[27\] VGND VGND VPWR VPWR net1774 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold544 CPU.registerFile\[26\]\[18\] VGND VGND VPWR VPWR net1785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 CPU.registerFile\[3\]\[21\] VGND VGND VPWR VPWR net1796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 CPU.registerFile\[12\]\[31\] VGND VGND VPWR VPWR net1807 sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 CPU.registerFile\[20\]\[2\] VGND VGND VPWR VPWR net1818 sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 CPU.registerFile\[26\]\[25\] VGND VGND VPWR VPWR net1829 sky130_fd_sc_hd__dlygate4sd3_1
X_09954_ _05509_ net1614 _05559_ VGND VGND VPWR VPWR _05569_ sky130_fd_sc_hd__mux2_1
Xhold599 CPU.registerFile\[14\]\[15\] VGND VGND VPWR VPWR net1840 sky130_fd_sc_hd__dlygate4sd3_1
X_08905_ _04484_ _04624_ VGND VGND VPWR VPWR _04625_ sky130_fd_sc_hd__nor2_1
X_09885_ _05524_ net2241 _05512_ VGND VGND VPWR VPWR _05525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1200 mapped_spi_flash.rcv_data\[9\] VGND VGND VPWR VPWR net2441 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1211 CPU.aluReg\[31\] VGND VGND VPWR VPWR net2452 sky130_fd_sc_hd__dlygate4sd3_1
X_08836_ CPU.aluIn1\[13\] CPU.aluIn1\[12\] _04494_ VGND VGND VPWR VPWR _04556_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_146_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1222 CPU.registerFile\[17\]\[8\] VGND VGND VPWR VPWR net2463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1233 CPU.aluReg\[29\] VGND VGND VPWR VPWR net2474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1244 mapped_spi_ram.rcv_data\[8\] VGND VGND VPWR VPWR net2485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1255 CPU.aluIn1\[8\] VGND VGND VPWR VPWR net2496 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1266 CPU.registerFile\[7\]\[21\] VGND VGND VPWR VPWR net2507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1277 CPU.registerFile\[6\]\[12\] VGND VGND VPWR VPWR net2518 sky130_fd_sc_hd__dlygate4sd3_1
X_08767_ CPU.Jimm\[13\] CPU.Jimm\[12\] VGND VGND VPWR VPWR _04487_ sky130_fd_sc_hd__nor2_4
Xhold1288 mapped_spi_flash.div_counter\[0\] VGND VGND VPWR VPWR net2529 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_406 _04659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14465__592 clknet_1_0__leaf__02662_ VGND VGND VPWR VPWR net624 sky130_fd_sc_hd__inv_2
Xhold1299 mapped_spi_flash.rbusy VGND VGND VPWR VPWR net2540 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_417 _02856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08698_ _04408_ _04416_ _04417_ VGND VGND VPWR VPWR _04418_ sky130_fd_sc_hd__o21a_1
XFILLER_0_95_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10660_ _00004_ _06014_ _06017_ VGND VGND VPWR VPWR _06018_ sky130_fd_sc_hd__nand3b_4
XTAP_TAPCELL_ROW_62_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09319_ _05026_ VGND VGND VPWR VPWR _05027_ sky130_fd_sc_hd__buf_6
XFILLER_0_35_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10591_ net1404 _05970_ VGND VGND VPWR VPWR _05977_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_11_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12330_ _06981_ VGND VGND VPWR VPWR _01420_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12261_ CPU.aluIn1\[14\] _06930_ _06927_ VGND VGND VPWR VPWR _06931_ sky130_fd_sc_hd__mux2_1
X_11212_ _05541_ net2136 _06310_ VGND VGND VPWR VPWR _06315_ sky130_fd_sc_hd__mux2_1
X_14630__740 clknet_1_1__leaf__02679_ VGND VGND VPWR VPWR net772 sky130_fd_sc_hd__inv_2
XFILLER_0_102_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput7 net7 VGND VGND VPWR VPWR spi_clk sky130_fd_sc_hd__clkbuf_4
X_12192_ CPU.aluIn1\[30\] _06877_ _06865_ VGND VGND VPWR VPWR _06878_ sky130_fd_sc_hd__mux2_1
X_11143_ _06278_ VGND VGND VPWR VPWR _01942_ sky130_fd_sc_hd__clkbuf_1
X_15951_ _02759_ _03431_ _03433_ _03019_ VGND VGND VPWR VPWR _03434_ sky130_fd_sc_hd__a211o_1
X_11074_ _06241_ VGND VGND VPWR VPWR _01974_ sky130_fd_sc_hd__clkbuf_1
X_14548__667 clknet_1_1__leaf__02670_ VGND VGND VPWR VPWR net699 sky130_fd_sc_hd__inv_2
X_14969__1046 clknet_1_0__leaf__02712_ VGND VGND VPWR VPWR net1078 sky130_fd_sc_hd__inv_2
X_10025_ _05595_ VGND VGND VPWR VPWR _05607_ sky130_fd_sc_hd__buf_4
X_15882_ CPU.registerFile\[12\]\[14\] _03118_ VGND VGND VPWR VPWR _03367_ sky130_fd_sc_hd__or2_1
X_17621_ net810 _01909_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17552_ net741 _01840_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_11976_ _04933_ net1835 _06747_ VGND VGND VPWR VPWR _06756_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13715_ _07351_ _08133_ VGND VGND VPWR VPWR _08134_ sky130_fd_sc_hd__or2_1
XFILLER_0_156_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10927_ _06163_ VGND VGND VPWR VPWR _02043_ sky130_fd_sc_hd__clkbuf_1
X_17483_ net672 _01771_ VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dfxtp_1
X_14695_ clknet_1_1__leaf__02675_ VGND VGND VPWR VPWR _02685_ sky130_fd_sc_hd__buf_1
XFILLER_0_156_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13646_ _07818_ _08065_ _08066_ VGND VGND VPWR VPWR _08067_ sky130_fd_sc_hd__o21a_1
X_16434_ _02945_ _03900_ _03902_ _02864_ VGND VGND VPWR VPWR _03903_ sky130_fd_sc_hd__a211o_1
X_10858_ _06126_ VGND VGND VPWR VPWR _02075_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16365_ CPU.registerFile\[9\]\[28\] _02802_ _02803_ VGND VGND VPWR VPWR _03836_ sky130_fd_sc_hd__o21a_1
X_13577_ _07646_ _07989_ _07992_ _07999_ VGND VGND VPWR VPWR _08000_ sky130_fd_sc_hd__a31o_1
XFILLER_0_125_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10789_ _05528_ net2045 _06081_ VGND VGND VPWR VPWR _06090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15316_ CPU.registerFile\[5\]\[0\] CPU.registerFile\[4\]\[0\] _02805_ VGND VGND VPWR
+ VPWR _02815_ sky130_fd_sc_hd__mux2_1
X_18104_ net167 _02384_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_14713__815 clknet_1_0__leaf__02687_ VGND VGND VPWR VPWR net847 sky130_fd_sc_hd__inv_2
X_12528_ _07086_ VGND VGND VPWR VPWR _01294_ sky130_fd_sc_hd__clkbuf_1
X_16296_ CPU.registerFile\[15\]\[26\] _02826_ _02770_ _03768_ VGND VGND VPWR VPWR
+ _03769_ sky130_fd_sc_hd__o211a_1
XFILLER_0_124_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14293__437 clknet_1_0__leaf__08462_ VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__inv_2
XFILLER_0_152_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18035_ net1208 _02315_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[29\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_113_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12459_ net1933 _05668_ _07049_ VGND VGND VPWR VPWR _07050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14129_ mapped_spi_ram.rcv_data\[23\] _04688_ _04690_ mapped_spi_flash.rcv_data\[23\]
+ VGND VGND VPWR VPWR _08394_ sky130_fd_sc_hd__a22o_4
XFILLER_0_94_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09670_ mapped_spi_flash.rcv_data\[27\] _04709_ _04643_ per_uart.rx_data\[3\] VGND
+ VGND VPWR VPWR _05362_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08621_ CPU.aluIn1\[20\] _04246_ VGND VGND VPWR VPWR _04341_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17819_ net1008 _02103_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08552_ CPU.mem_wdata\[7\] CPU.Bimm\[7\] net1295 VGND VGND VPWR VPWR _04272_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_124_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_141_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08483_ _04202_ VGND VGND VPWR VPWR _04203_ sky130_fd_sc_hd__buf_6
XFILLER_0_76_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09104_ _04196_ _04372_ CPU.instr\[2\] VGND VGND VPWR VPWR _04816_ sky130_fd_sc_hd__or3b_1
XFILLER_0_45_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_749 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09035_ _04356_ _04469_ _04733_ VGND VGND VPWR VPWR _04750_ sky130_fd_sc_hd__nor3_1
Xhold330 CPU.registerFile\[8\]\[26\] VGND VGND VPWR VPWR net1571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 CPU.registerFile\[8\]\[30\] VGND VGND VPWR VPWR net1582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 per_uart.uart0.tx_count16\[3\] VGND VGND VPWR VPWR net1593 sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 CPU.registerFile\[5\]\[11\] VGND VGND VPWR VPWR net1604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 CPU.registerFile\[4\]\[1\] VGND VGND VPWR VPWR net1615 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold385 CPU.registerFile\[6\]\[2\] VGND VGND VPWR VPWR net1626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 per_uart.d_in_uart\[1\] VGND VGND VPWR VPWR net1637 sky130_fd_sc_hd__dlygate4sd3_1
X_09937_ _05560_ VGND VGND VPWR VPWR _02477_ sky130_fd_sc_hd__clkbuf_1
X_09868_ _05513_ VGND VGND VPWR VPWR _02499_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1030 CPU.registerFile\[31\]\[0\] VGND VGND VPWR VPWR net2271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1041 CPU.registerFile\[19\]\[7\] VGND VGND VPWR VPWR net2282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1052 CPU.registerFile\[15\]\[7\] VGND VGND VPWR VPWR net2293 sky130_fd_sc_hd__dlygate4sd3_1
X_08819_ CPU.aluIn1\[6\] CPU.Bimm\[6\] VGND VGND VPWR VPWR _04539_ sky130_fd_sc_hd__and2_1
Xhold1063 CPU.registerFile\[27\]\[3\] VGND VGND VPWR VPWR net2304 sky130_fd_sc_hd__dlygate4sd3_1
X_09799_ _05470_ VGND VGND VPWR VPWR _02525_ sky130_fd_sc_hd__clkbuf_1
Xhold1074 CPU.registerFile\[28\]\[8\] VGND VGND VPWR VPWR net2315 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1085 CPU.registerFile\[22\]\[18\] VGND VGND VPWR VPWR net2326 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_203 _07841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11830_ net2144 _05677_ _06675_ VGND VGND VPWR VPWR _06679_ sky130_fd_sc_hd__mux2_1
Xhold1096 CPU.registerFile\[28\]\[4\] VGND VGND VPWR VPWR net2337 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_214 _07999_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_225 clknet_1_0__leaf__02720_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_236 _02873_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_247 _03330_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11761_ _06642_ VGND VGND VPWR VPWR _01685_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_258 _05050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_269 _05448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13500_ CPU.registerFile\[23\]\[18\] _07362_ _07619_ CPU.registerFile\[19\]\[18\]
+ _07924_ VGND VGND VPWR VPWR _07925_ sky130_fd_sc_hd__o221a_1
X_10712_ _06049_ VGND VGND VPWR VPWR _02144_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11692_ mapped_spi_ram.rcv_data\[14\] _06588_ VGND VGND VPWR VPWR _06599_ sky130_fd_sc_hd__or2_1
X_13431_ CPU.registerFile\[30\]\[15\] CPU.registerFile\[26\]\[15\] _07352_ VGND VGND
+ VPWR VPWR _07859_ sky130_fd_sc_hd__mux2_1
X_10643_ net1500 _05996_ _06005_ _06006_ VGND VGND VPWR VPWR _02169_ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16150_ _02926_ _03626_ _03627_ VGND VGND VPWR VPWR _03628_ sky130_fd_sc_hd__o21a_1
X_13362_ CPU.registerFile\[28\]\[13\] CPU.registerFile\[24\]\[13\] _07292_ VGND VGND
+ VPWR VPWR _07792_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10574_ _05962_ _05965_ VGND VGND VPWR VPWR _05966_ sky130_fd_sc_hd__or2b_1
X_15101_ _07189_ _02737_ _02727_ VGND VGND VPWR VPWR _02280_ sky130_fd_sc_hd__a21oi_1
Xrebuffer8 net1250 VGND VGND VPWR VPWR net1249 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12313_ CPU.aluReg\[2\] CPU.aluReg\[0\] _06870_ VGND VGND VPWR VPWR _06970_ sky130_fd_sc_hd__mux2_1
X_16081_ CPU.registerFile\[30\]\[19\] _05050_ _02923_ _03560_ VGND VGND VPWR VPWR
+ _03561_ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13293_ CPU.registerFile\[29\]\[11\] _07403_ _07404_ CPU.registerFile\[25\]\[11\]
+ _07250_ VGND VGND VPWR VPWR _07725_ sky130_fd_sc_hd__o221a_1
X_12244_ CPU.aluReg\[18\] _06917_ _06891_ VGND VGND VPWR VPWR _06918_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12175_ _06859_ VGND VGND VPWR VPWR _06865_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_75_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11126_ _06269_ VGND VGND VPWR VPWR _01950_ sky130_fd_sc_hd__clkbuf_1
X_16983_ clknet_leaf_21_clk _01309_ VGND VGND VPWR VPWR CPU.rs2\[14\] sky130_fd_sc_hd__dfxtp_1
X_11057_ _06232_ VGND VGND VPWR VPWR _01982_ sky130_fd_sc_hd__clkbuf_1
X_15934_ CPU.registerFile\[25\]\[15\] CPU.registerFile\[29\]\[15\] _02851_ VGND VGND
+ VPWR VPWR _03418_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14481__607 clknet_1_0__leaf__02663_ VGND VGND VPWR VPWR net639 sky130_fd_sc_hd__inv_2
X_10008_ _05598_ VGND VGND VPWR VPWR _02412_ sky130_fd_sc_hd__clkbuf_1
X_15865_ CPU.registerFile\[7\]\[13\] _03317_ VGND VGND VPWR VPWR _03351_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17604_ net793 _01892_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_15796_ CPU.registerFile\[7\]\[11\] _05092_ VGND VGND VPWR VPWR _03284_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_35_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_646 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17535_ net724 _01823_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11959_ _06746_ VGND VGND VPWR VPWR _06747_ sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_103_Left_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17466_ net655 _01754_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13629_ CPU.registerFile\[6\]\[22\] CPU.registerFile\[7\]\[22\] _07641_ VGND VGND
+ VPWR VPWR _08050_ sky130_fd_sc_hd__mux2_1
X_16417_ CPU.registerFile\[25\]\[29\] CPU.registerFile\[29\]\[29\] _03254_ VGND VGND
+ VPWR VPWR _03887_ sky130_fd_sc_hd__mux2_1
X_17397_ net586 _01685_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_14301__444 clknet_1_1__leaf__08463_ VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__inv_2
XFILLER_0_6_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16348_ CPU.registerFile\[28\]\[27\] _02772_ VGND VGND VPWR VPWR _03820_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16279_ CPU.registerFile\[16\]\[25\] CPU.registerFile\[18\]\[25\] _05440_ VGND VGND
+ VPWR VPWR _03753_ sky130_fd_sc_hd__mux2_1
X_18018_ net1191 _02298_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_112_Left_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09722_ _04873_ _05411_ VGND VGND VPWR VPWR _05412_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_126_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09653_ CPU.PC\[3\] CPU.PC\[2\] CPU.PC\[4\] VGND VGND VPWR VPWR _05346_ sky130_fd_sc_hd__a21oi_1
X_08604_ _04323_ _04319_ _04321_ VGND VGND VPWR VPWR _04324_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09584_ mapped_spi_flash.rcv_data\[30\] _04784_ _05278_ VGND VGND VPWR VPWR _05279_
+ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_121_Left_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_118_Right_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08535_ CPU.rs2\[15\] _04200_ _04205_ VGND VGND VPWR VPWR _04255_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_526 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14577__693 clknet_1_0__leaf__02673_ VGND VGND VPWR VPWR net725 sky130_fd_sc_hd__inv_2
X_14968__1045 clknet_1_0__leaf__02712_ VGND VGND VPWR VPWR net1077 sky130_fd_sc_hd__inv_2
XFILLER_0_122_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09018_ _04469_ _04733_ _04356_ VGND VGND VPWR VPWR _04734_ sky130_fd_sc_hd__o21a_1
X_10290_ _05764_ VGND VGND VPWR VPWR _02296_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold160 mapped_spi_flash.cmd_addr\[18\] VGND VGND VPWR VPWR net1401 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 mapped_spi_ram.rcv_data\[26\] VGND VGND VPWR VPWR net1412 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold182 per_uart.uart0.enable16_counter\[4\] VGND VGND VPWR VPWR net1423 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 mapped_spi_ram.rcv_data\[24\] VGND VGND VPWR VPWR net1434 sky130_fd_sc_hd__dlygate4sd3_1
X_14742__841 clknet_1_0__leaf__02690_ VGND VGND VPWR VPWR net873 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_70_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12931_ CPU.registerFile\[6\]\[2\] CPU.registerFile\[7\]\[2\] _07371_ VGND VGND VPWR
+ VPWR _07372_ sky130_fd_sc_hd__mux2_1
X_16502__171 clknet_1_1__leaf__03962_ VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__inv_2
X_15650_ CPU.registerFile\[6\]\[7\] _03057_ _03140_ _03141_ VGND VGND VPWR VPWR _03142_
+ sky130_fd_sc_hd__o211a_1
X_12862_ _07304_ VGND VGND VPWR VPWR _07305_ sky130_fd_sc_hd__buf_4
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11813_ _06669_ VGND VGND VPWR VPWR _01660_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15581_ CPU.registerFile\[18\]\[5\] _02832_ _02835_ CPU.registerFile\[19\]\[5\] _03074_
+ VGND VGND VPWR VPWR _03075_ sky130_fd_sc_hd__o221a_1
XFILLER_0_68_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12793_ _07235_ VGND VGND VPWR VPWR _07236_ sky130_fd_sc_hd__buf_4
XFILLER_0_139_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17320_ net509 _01608_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11744_ _06571_ _06631_ VGND VGND VPWR VPWR _06632_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17251_ net441 _01539_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11675_ net1448 _06575_ _06589_ _06581_ VGND VGND VPWR VPWR _01717_ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13414_ CPU.registerFile\[6\]\[15\] CPU.registerFile\[7\]\[15\] _07263_ VGND VGND
+ VPWR VPWR _07842_ sky130_fd_sc_hd__mux2_1
X_16202_ _03227_ _03672_ _03673_ _03228_ _03677_ VGND VGND VPWR VPWR _03678_ sky130_fd_sc_hd__a221o_1
XFILLER_0_126_559 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17182_ clknet_leaf_14_clk _01470_ VGND VGND VPWR VPWR CPU.Jimm\[12\] sky130_fd_sc_hd__dfxtp_1
X_10626_ net2064 _05996_ _05997_ _05993_ VGND VGND VPWR VPWR _02177_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16133_ _02911_ _03608_ _03610_ _03245_ VGND VGND VPWR VPWR _03611_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_77_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13345_ _07370_ _07774_ VGND VGND VPWR VPWR _07775_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_77_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10557_ _05945_ _05953_ VGND VGND VPWR VPWR _05954_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16064_ _02949_ _03540_ _03543_ VGND VGND VPWR VPWR _03544_ sky130_fd_sc_hd__or3_4
X_13276_ CPU.registerFile\[23\]\[11\] _07362_ _07619_ CPU.registerFile\[19\]\[11\]
+ _07707_ VGND VGND VPWR VPWR _07708_ sky130_fd_sc_hd__o221a_2
X_10488_ net1400 _05892_ _05897_ _05885_ VGND VGND VPWR VPWR _02215_ sky130_fd_sc_hd__o211a_1
X_12227_ CPU.aluReg\[22\] _06904_ _06891_ VGND VGND VPWR VPWR _06905_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_90_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14825__916 clknet_1_1__leaf__02698_ VGND VGND VPWR VPWR net948 sky130_fd_sc_hd__inv_2
X_12158_ _05426_ net2410 _06818_ VGND VGND VPWR VPWR _06852_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11109_ _06260_ VGND VGND VPWR VPWR _01958_ sky130_fd_sc_hd__clkbuf_1
X_16966_ net261 _01292_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_12089_ _06815_ VGND VGND VPWR VPWR _01529_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_108_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15917_ _03399_ _03400_ _02856_ VGND VGND VPWR VPWR _03401_ sky130_fd_sc_hd__mux2_1
X_16897_ _04148_ _04174_ VGND VGND VPWR VPWR _04175_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15848_ CPU.registerFile\[12\]\[13\] _03118_ VGND VGND VPWR VPWR _03334_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_88_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_121_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15779_ CPU.registerFile\[8\]\[11\] _02763_ _03117_ _03266_ VGND VGND VPWR VPWR _03267_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17518_ net707 _01806_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14871__958 clknet_1_1__leaf__02702_ VGND VGND VPWR VPWR net990 sky130_fd_sc_hd__inv_2
XFILLER_0_90_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17449_ net638 _01737_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09705_ net1293 _04304_ VGND VGND VPWR VPWR _05396_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09636_ CPU.cycles\[5\] _04502_ VGND VGND VPWR VPWR _05330_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09567_ _05262_ _04424_ VGND VGND VPWR VPWR _05263_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_616 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08518_ CPU.aluIn1\[23\] _04237_ VGND VGND VPWR VPWR _04238_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_26_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09498_ _04921_ _05196_ VGND VGND VPWR VPWR _05197_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_156_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11460_ _05516_ net2033 _06444_ VGND VGND VPWR VPWR _06447_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_816 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10411_ mapped_spi_flash.cmd_addr\[26\] _05825_ _05827_ mapped_spi_flash.cmd_addr\[27\]
+ VGND VGND VPWR VPWR _05837_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_59_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11391_ _06410_ VGND VGND VPWR VPWR _01826_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13130_ CPU.mem_wdata\[6\] _07229_ _07566_ _07135_ VGND VGND VPWR VPWR _01301_ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10342_ _05792_ VGND VGND VPWR VPWR _02257_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13061_ _07322_ _07498_ VGND VGND VPWR VPWR _07499_ sky130_fd_sc_hd__or2_1
X_10273_ _05755_ VGND VGND VPWR VPWR _02304_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_72_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12012_ _05306_ net2486 _06769_ VGND VGND VPWR VPWR _06775_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16820_ net1593 VGND VGND VPWR VPWR _04123_ sky130_fd_sc_hd__inv_2
X_14330__470 clknet_1_0__leaf__08466_ VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__inv_2
X_16751_ _04001_ _05101_ VGND VGND VPWR VPWR _04069_ sky130_fd_sc_hd__nand2_1
X_15702_ CPU.registerFile\[14\]\[9\] CPU.registerFile\[10\]\[9\] _02849_ VGND VGND
+ VPWR VPWR _03192_ sky130_fd_sc_hd__mux2_1
X_12914_ _07271_ _07338_ _07342_ _07355_ _07306_ VGND VGND VPWR VPWR _07356_ sky130_fd_sc_hd__o311a_1
X_13894_ CPU.registerFile\[1\]\[30\] _07255_ _08306_ _07318_ VGND VGND VPWR VPWR _08307_
+ sky130_fd_sc_hd__a22o_1
X_16682_ _03991_ net1549 VGND VGND VPWR VPWR _04010_ sky130_fd_sc_hd__nand2_1
X_15633_ _02779_ VGND VGND VPWR VPWR _03125_ sky130_fd_sc_hd__clkbuf_4
X_12845_ _07252_ VGND VGND VPWR VPWR _07288_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_103_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18352_ clknet_leaf_6_clk _02632_ VGND VGND VPWR VPWR per_uart.uart0.rx_bitcount\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15564_ CPU.registerFile\[7\]\[5\] _05092_ VGND VGND VPWR VPWR _03058_ sky130_fd_sc_hd__or2_1
X_14593__708 clknet_1_1__leaf__02674_ VGND VGND VPWR VPWR net740 sky130_fd_sc_hd__inv_2
XFILLER_0_139_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17303_ net492 _01591_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11727_ net8 net22 _06617_ net1309 _04589_ VGND VGND VPWR VPWR _06619_ sky130_fd_sc_hd__a41o_1
X_18283_ net116 _02563_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15495_ _02827_ _02989_ _02990_ VGND VGND VPWR VPWR _02991_ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17234_ net424 _01522_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11658_ net1407 _06577_ VGND VGND VPWR VPWR _06580_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10609_ net1484 _05983_ _05987_ _05980_ VGND VGND VPWR VPWR _02184_ sky130_fd_sc_hd__o211a_1
X_17165_ net389 _01453_ VGND VGND VPWR VPWR CPU.aluReg\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11589_ _06512_ _05929_ VGND VGND VPWR VPWR _06531_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold907 CPU.registerFile\[11\]\[27\] VGND VGND VPWR VPWR net2148 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__08430_ _08430_ VGND VGND VPWR VPWR clknet_0__08430_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16116_ CPU.registerFile\[30\]\[20\] _05050_ _02923_ _03594_ VGND VGND VPWR VPWR
+ _03595_ sky130_fd_sc_hd__o211a_1
X_13328_ CPU.registerFile\[30\]\[12\] CPU.registerFile\[26\]\[12\] _07297_ VGND VGND
+ VPWR VPWR _07759_ sky130_fd_sc_hd__mux2_1
Xhold918 CPU.registerFile\[23\]\[23\] VGND VGND VPWR VPWR net2159 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12771__220 clknet_1_0__leaf__07225_ VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__inv_2
XFILLER_0_122_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17096_ net354 _01418_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[26\] sky130_fd_sc_hd__dfxtp_1
Xhold929 CPU.registerFile\[20\]\[29\] VGND VGND VPWR VPWR net2170 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__02754_ clknet_0__02754_ VGND VGND VPWR VPWR clknet_1_1__leaf__02754_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_40_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__08361_ _08361_ VGND VGND VPWR VPWR clknet_0__08361_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_150_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13259_ CPU.registerFile\[30\]\[10\] CPU.registerFile\[26\]\[10\] _04937_ VGND VGND
+ VPWR VPWR _07692_ sky130_fd_sc_hd__mux2_1
X_16047_ _05010_ _03524_ _03527_ VGND VGND VPWR VPWR _03528_ sky130_fd_sc_hd__or3_2
XFILLER_0_20_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14413__545 clknet_1_1__leaf__02657_ VGND VGND VPWR VPWR net577 sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__02685_ clknet_0__02685_ VGND VGND VPWR VPWR clknet_1_1__leaf__02685_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17998_ clknet_leaf_7_clk _02282_ VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_16949_ net244 _01275_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_14967__1044 clknet_1_1__leaf__02712_ VGND VGND VPWR VPWR net1076 sky130_fd_sc_hd__inv_2
XFILLER_0_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09421_ CPU.PC\[14\] _04846_ VGND VGND VPWR VPWR _05124_ sky130_fd_sc_hd__xor2_1
XFILLER_0_94_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09352_ _04253_ _04683_ VGND VGND VPWR VPWR _05058_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09283_ _04342_ _04699_ _04808_ CPU.aluReg\[20\] _04991_ VGND VGND VPWR VPWR _04992_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload80 clknet_1_0__leaf__02653_ VGND VGND VPWR VPWR clkload80/X sky130_fd_sc_hd__clkbuf_8
Xclkload91 clknet_1_1__leaf__08468_ VGND VGND VPWR VPWR clkload91/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_30_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14689__794 clknet_1_1__leaf__02684_ VGND VGND VPWR VPWR net826 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_54_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14388__522 clknet_1_1__leaf__02655_ VGND VGND VPWR VPWR net554 sky130_fd_sc_hd__inv_2
X_08998_ _04715_ VGND VGND VPWR VPWR _02579_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_149_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10960_ _06181_ VGND VGND VPWR VPWR _02028_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09619_ _04624_ _04621_ VGND VGND VPWR VPWR _05313_ sky130_fd_sc_hd__nand2_1
X_10891_ net1550 _05673_ _06143_ VGND VGND VPWR VPWR _06145_ sky130_fd_sc_hd__mux2_1
X_12630_ net1501 _07138_ VGND VGND VPWR VPWR _00041_ sky130_fd_sc_hd__xor2_1
XFILLER_0_127_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14854__942 clknet_1_0__leaf__02701_ VGND VGND VPWR VPWR net974 sky130_fd_sc_hd__inv_2
X_12561_ _07103_ VGND VGND VPWR VPWR _01278_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11512_ _06030_ _06477_ VGND VGND VPWR VPWR _01772_ sky130_fd_sc_hd__nor2_1
X_15280_ _05069_ VGND VGND VPWR VPWR _02779_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_25_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12492_ net1947 _05704_ _07060_ VGND VGND VPWR VPWR _07067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11443_ _05499_ CPU.registerFile\[25\]\[27\] _06433_ VGND VGND VPWR VPWR _06438_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14162_ CPU.Iimm\[4\] _07232_ _08413_ VGND VGND VPWR VPWR _08418_ sky130_fd_sc_hd__mux2_1
X_11374_ _06401_ VGND VGND VPWR VPWR _01834_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13113_ CPU.registerFile\[13\]\[6\] _07382_ _07549_ VGND VGND VPWR VPWR _07550_ sky130_fd_sc_hd__o21a_1
XFILLER_0_150_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10325_ _05783_ VGND VGND VPWR VPWR _02265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14093_ _08373_ VGND VGND VPWR VPWR _01457_ sky130_fd_sc_hd__clkbuf_1
X_13044_ _05308_ VGND VGND VPWR VPWR _07483_ sky130_fd_sc_hd__buf_4
X_17921_ net1110 _02205_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[1\] sky130_fd_sc_hd__dfxtp_1
X_10256_ _05746_ VGND VGND VPWR VPWR _02312_ sky130_fd_sc_hd__clkbuf_1
X_17852_ net1041 _02136_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_10187_ net2368 _05700_ _05692_ VGND VGND VPWR VPWR _05701_ sky130_fd_sc_hd__mux2_1
X_16803_ net1537 VGND VGND VPWR VPWR _02604_ sky130_fd_sc_hd__clkbuf_1
X_17783_ net972 _02067_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_14995_ clknet_1_1__leaf__02708_ VGND VGND VPWR VPWR _02715_ sky130_fd_sc_hd__buf_1
X_16734_ _04050_ _04051_ _04053_ _04054_ VGND VGND VPWR VPWR _04055_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16665_ _03995_ _05396_ _07123_ VGND VGND VPWR VPWR _03996_ sky130_fd_sc_hd__o21ai_1
X_13877_ _07296_ _08290_ VGND VGND VPWR VPWR _08291_ sky130_fd_sc_hd__or2_1
X_15616_ _02827_ _03107_ _03108_ VGND VGND VPWR VPWR _03109_ sky130_fd_sc_hd__o21ai_1
X_12828_ _05232_ VGND VGND VPWR VPWR _07271_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_57_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18335_ clknet_leaf_9_clk _02615_ VGND VGND VPWR VPWR per_uart.uart0.txd_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_15547_ CPU.registerFile\[15\]\[5\] CPU.registerFile\[11\]\[5\] _02773_ VGND VGND
+ VPWR VPWR _03041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12759_ clknet_1_1__leaf__07223_ VGND VGND VPWR VPWR _07224_ sky130_fd_sc_hd__buf_1
XFILLER_0_44_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18266_ clknet_leaf_1_clk _02546_ VGND VGND VPWR VPWR per_uart.uart0.rxd_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15478_ CPU.registerFile\[25\]\[3\] _02943_ _02860_ VGND VGND VPWR VPWR _02974_ sky130_fd_sc_hd__o21a_1
XFILLER_0_112_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17217_ net407 _01505_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_14429_ clknet_1_1__leaf__02653_ VGND VGND VPWR VPWR _02659_ sky130_fd_sc_hd__buf_1
X_18197_ net228 _02477_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17148_ net372 _01436_ VGND VGND VPWR VPWR CPU.aluReg\[12\] sky130_fd_sc_hd__dfxtp_1
Xhold704 CPU.registerFile\[18\]\[3\] VGND VGND VPWR VPWR net1945 sky130_fd_sc_hd__dlygate4sd3_1
Xhold715 CPU.registerFile\[13\]\[3\] VGND VGND VPWR VPWR net1956 sky130_fd_sc_hd__dlygate4sd3_1
Xhold726 CPU.registerFile\[1\]\[11\] VGND VGND VPWR VPWR net1967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold737 CPU.registerFile\[1\]\[6\] VGND VGND VPWR VPWR net1978 sky130_fd_sc_hd__dlygate4sd3_1
X_09970_ _05577_ VGND VGND VPWR VPWR _02461_ sky130_fd_sc_hd__clkbuf_1
Xhold748 CPU.registerFile\[22\]\[4\] VGND VGND VPWR VPWR net1989 sky130_fd_sc_hd__dlygate4sd3_1
Xhold759 CPU.registerFile\[28\]\[18\] VGND VGND VPWR VPWR net2000 sky130_fd_sc_hd__dlygate4sd3_1
X_17079_ net337 _01401_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08921_ _04616_ _04615_ _04612_ _04640_ VGND VGND VPWR VPWR _04641_ sky130_fd_sc_hd__and4_1
XFILLER_0_0_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__02668_ clknet_0__02668_ VGND VGND VPWR VPWR clknet_1_1__leaf__02668_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08852_ CPU.aluIn1\[20\] _04495_ VGND VGND VPWR VPWR _04572_ sky130_fd_sc_hd__nand2_1
Xclkbuf_0__02699_ _02699_ VGND VGND VPWR VPWR clknet_0__02699_ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_0__07226_ _07226_ VGND VGND VPWR VPWR clknet_0__07226_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_137_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08783_ _04502_ VGND VGND VPWR VPWR _04503_ sky130_fd_sc_hd__clkbuf_4
X_15238__147 clknet_1_0__leaf__02754_ VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14012__292 clknet_1_1__leaf__08361_ VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__inv_2
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09404_ _04717_ _05094_ _05098_ _05107_ VGND VGND VPWR VPWR _05108_ sky130_fd_sc_hd__a211o_4
XFILLER_0_94_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09335_ _04902_ _05041_ VGND VGND VPWR VPWR _05042_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09266_ CPU.PC\[21\] _04928_ VGND VGND VPWR VPWR _04976_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09197_ CPU.PC\[22\] _04821_ _04908_ VGND VGND VPWR VPWR _04909_ sky130_fd_sc_hd__o21a_1
XFILLER_0_90_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10110_ _05652_ VGND VGND VPWR VPWR _02364_ sky130_fd_sc_hd__clkbuf_1
X_11090_ _06249_ VGND VGND VPWR VPWR _01966_ sky130_fd_sc_hd__clkbuf_1
X_10041_ _05615_ VGND VGND VPWR VPWR _02396_ sky130_fd_sc_hd__clkbuf_1
Xhold75 mapped_spi_flash.rcv_data\[30\] VGND VGND VPWR VPWR net1316 sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ CPU.registerFile\[21\]\[27\] _07244_ _07429_ CPU.registerFile\[17\]\[27\]
+ _07349_ VGND VGND VPWR VPWR _08216_ sky130_fd_sc_hd__o221a_1
Xhold86 mapped_spi_ram.cmd_addr\[29\] VGND VGND VPWR VPWR net1327 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 _02165_ VGND VGND VPWR VPWR net1338 sky130_fd_sc_hd__dlygate4sd3_1
X_11992_ _06764_ VGND VGND VPWR VPWR _01576_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10943_ net1581 _05725_ _06165_ VGND VGND VPWR VPWR _06172_ sky130_fd_sc_hd__mux2_1
X_13731_ _08146_ _08147_ _08148_ _04814_ _07272_ VGND VGND VPWR VPWR _08149_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_67_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16450_ _02848_ _03914_ _03918_ _02843_ VGND VGND VPWR VPWR _03919_ sky130_fd_sc_hd__a211o_1
XFILLER_0_97_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10874_ net2070 _05725_ _06128_ VGND VGND VPWR VPWR _06135_ sky130_fd_sc_hd__mux2_1
X_13662_ _07987_ _04987_ VGND VGND VPWR VPWR _08082_ sky130_fd_sc_hd__nor2_1
X_14442__571 clknet_1_1__leaf__02660_ VGND VGND VPWR VPWR net603 sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__02688_ clknet_0__02688_ VGND VGND VPWR VPWR clknet_1_0__leaf__02688_
+ sky130_fd_sc_hd__clkbuf_16
X_15401_ _02896_ _02897_ _02898_ VGND VGND VPWR VPWR _02899_ sky130_fd_sc_hd__mux2_1
X_12613_ net21 _06493_ _04192_ VGND VGND VPWR VPWR _07130_ sky130_fd_sc_hd__and3b_1
X_16381_ _08404_ _03850_ _03851_ VGND VGND VPWR VPWR _03852_ sky130_fd_sc_hd__a21o_1
X_13593_ _07394_ _08000_ _08014_ _08015_ VGND VGND VPWR VPWR _08016_ sky130_fd_sc_hd__a211o_1
XFILLER_0_155_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18120_ net183 _02400_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12544_ _07094_ VGND VGND VPWR VPWR _01286_ sky130_fd_sc_hd__clkbuf_1
X_15332_ _04620_ _05048_ VGND VGND VPWR VPWR _02831_ sky130_fd_sc_hd__nand2_2
XFILLER_0_54_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18051_ net1224 _02331_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_12475_ net1844 _05687_ _07049_ VGND VGND VPWR VPWR _07058_ sky130_fd_sc_hd__mux2_1
X_15263_ CPU.registerFile\[14\]\[0\] CPU.registerFile\[10\]\[0\] _02761_ VGND VGND
+ VPWR VPWR _02762_ sky130_fd_sc_hd__mux2_1
X_14966__1043 clknet_1_1__leaf__02712_ VGND VGND VPWR VPWR net1075 sky130_fd_sc_hd__inv_2
X_17002_ clknet_leaf_12_clk _00000_ VGND VGND VPWR VPWR CPU.state\[1\] sky130_fd_sc_hd__dfxtp_1
X_11426_ _06428_ VGND VGND VPWR VPWR _01809_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_6 _02800_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14145_ _05384_ VGND VGND VPWR VPWR _08407_ sky130_fd_sc_hd__clkbuf_4
X_11357_ _06391_ VGND VGND VPWR VPWR _01841_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10308_ _05773_ VGND VGND VPWR VPWR _02287_ sky130_fd_sc_hd__clkbuf_1
X_14076_ clknet_1_1__leaf__08363_ VGND VGND VPWR VPWR _08368_ sky130_fd_sc_hd__buf_1
X_11288_ CPU.registerFile\[9\]\[3\] _05729_ _06346_ VGND VGND VPWR VPWR _06355_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17904_ net1093 net1415 VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[22\] sky130_fd_sc_hd__dfxtp_1
X_13027_ CPU.registerFile\[16\]\[4\] CPU.registerFile\[20\]\[4\] _07339_ VGND VGND
+ VPWR VPWR _07466_ sky130_fd_sc_hd__mux2_1
X_10239_ net2208 _05735_ _05670_ VGND VGND VPWR VPWR _05736_ sky130_fd_sc_hd__mux2_1
X_17835_ net1024 _02119_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_17766_ net955 _02050_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[20\] sky130_fd_sc_hd__dfxtp_1
Xrebuffer18 net1260 VGND VGND VPWR VPWR net1259 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer29 net1271 VGND VGND VPWR VPWR net1270 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_16_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14525__646 clknet_1_0__leaf__02668_ VGND VGND VPWR VPWR net678 sky130_fd_sc_hd__inv_2
X_16717_ _04027_ _04039_ _05195_ VGND VGND VPWR VPWR _04040_ sky130_fd_sc_hd__a21o_1
X_13929_ CPU.registerFile\[15\]\[31\] _07236_ _07239_ CPU.registerFile\[11\]\[31\]
+ _07820_ VGND VGND VPWR VPWR _08341_ sky130_fd_sc_hd__o221a_1
X_17697_ net886 _01985_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09120_ CPU.Jimm\[19\] _04829_ _04831_ VGND VGND VPWR VPWR _04832_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18318_ clknet_leaf_15_clk _02598_ VGND VGND VPWR VPWR CPU.PC\[18\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_33_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09051_ _04733_ _04764_ VGND VGND VPWR VPWR _04765_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18249_ net90 _02529_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold501 CPU.registerFile\[26\]\[0\] VGND VGND VPWR VPWR net1742 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold512 CPU.registerFile\[3\]\[16\] VGND VGND VPWR VPWR net1753 sky130_fd_sc_hd__dlygate4sd3_1
X_14571__688 clknet_1_0__leaf__02672_ VGND VGND VPWR VPWR net720 sky130_fd_sc_hd__inv_2
Xhold523 CPU.registerFile\[12\]\[26\] VGND VGND VPWR VPWR net1764 sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 CPU.registerFile\[5\]\[14\] VGND VGND VPWR VPWR net1775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 CPU.registerFile\[29\]\[25\] VGND VGND VPWR VPWR net1786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 per_uart.uart0.rxd_reg\[6\] VGND VGND VPWR VPWR net1797 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold567 CPU.registerFile\[2\]\[4\] VGND VGND VPWR VPWR net1808 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold578 per_uart.d_in_uart\[4\] VGND VGND VPWR VPWR net1819 sky130_fd_sc_hd__dlygate4sd3_1
Xhold589 CPU.registerFile\[3\]\[9\] VGND VGND VPWR VPWR net1830 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ _05568_ VGND VGND VPWR VPWR _02469_ sky130_fd_sc_hd__clkbuf_1
X_08904_ _04524_ _04623_ VGND VGND VPWR VPWR _04624_ sky130_fd_sc_hd__nand2_2
X_09884_ _05108_ VGND VGND VPWR VPWR _05524_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_148_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1201 CPU.registerFile\[27\]\[19\] VGND VGND VPWR VPWR net2442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1212 CPU.registerFile\[9\]\[28\] VGND VGND VPWR VPWR net2453 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08835_ CPU.aluIn1\[14\] _04494_ VGND VGND VPWR VPWR _04555_ sky130_fd_sc_hd__xnor2_2
Xhold1223 CPU.registerFile\[25\]\[7\] VGND VGND VPWR VPWR net2464 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1234 CPU.registerFile\[25\]\[21\] VGND VGND VPWR VPWR net2475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1245 CPU.registerFile\[12\]\[6\] VGND VGND VPWR VPWR net2486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1256 CPU.aluIn1\[29\] VGND VGND VPWR VPWR net2497 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1267 CPU.registerFile\[7\]\[6\] VGND VGND VPWR VPWR net2508 sky130_fd_sc_hd__dlygate4sd3_1
X_08766_ _04374_ _04481_ _04482_ _04485_ VGND VGND VPWR VPWR _04486_ sky130_fd_sc_hd__a31o_1
Xhold1278 CPU.registerFile\[4\]\[15\] VGND VGND VPWR VPWR net2519 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1289 CPU.registerFile\[13\]\[6\] VGND VGND VPWR VPWR net2530 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_407 _04659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_418 _02856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08697_ _04305_ _04287_ VGND VGND VPWR VPWR _04417_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_49_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09318_ _05021_ _05012_ _05011_ _05025_ VGND VGND VPWR VPWR _05026_ sky130_fd_sc_hd__or4b_4
XTAP_TAPCELL_ROW_62_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10590_ net1404 _05968_ _05976_ _05936_ VGND VGND VPWR VPWR _02192_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_11_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_149_Left_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09249_ _04959_ VGND VGND VPWR VPWR _02572_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12260_ CPU.aluReg\[15\] CPU.aluReg\[13\] _06906_ VGND VGND VPWR VPWR _06930_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11211_ _06314_ VGND VGND VPWR VPWR _01910_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12191_ CPU.aluReg\[31\] CPU.aluReg\[29\] _06871_ VGND VGND VPWR VPWR _06877_ sky130_fd_sc_hd__mux2_1
Xoutput8 net8 VGND VGND VPWR VPWR spi_clk_ram sky130_fd_sc_hd__clkbuf_4
Xoutput10 net10 VGND VGND VPWR VPWR spi_cs_n_ram sky130_fd_sc_hd__buf_2
X_11142_ net2431 _05719_ _06274_ VGND VGND VPWR VPWR _06278_ sky130_fd_sc_hd__mux2_1
X_15950_ CPU.registerFile\[8\]\[16\] _02789_ _03117_ _03432_ VGND VGND VPWR VPWR _03433_
+ sky130_fd_sc_hd__o211a_1
X_11073_ net2460 _05719_ _06237_ VGND VGND VPWR VPWR _06241_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_158_Left_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10024_ _05606_ VGND VGND VPWR VPWR _02404_ sky130_fd_sc_hd__clkbuf_1
X_15881_ CPU.registerFile\[14\]\[14\] CPU.registerFile\[10\]\[14\] _03082_ VGND VGND
+ VPWR VPWR _03366_ sky130_fd_sc_hd__mux2_1
X_17620_ net809 _01908_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17551_ net740 _01839_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_11975_ _06755_ VGND VGND VPWR VPWR _01584_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13714_ CPU.registerFile\[30\]\[24\] CPU.registerFile\[26\]\[24\] _07297_ VGND VGND
+ VPWR VPWR _08133_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10926_ net1595 _05708_ _06154_ VGND VGND VPWR VPWR _06163_ sky130_fd_sc_hd__mux2_1
X_17482_ net671 net28 VGND VGND VPWR VPWR mapped_spi_flash.div_counter\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16578__50 clknet_1_1__leaf__03969_ VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__inv_2
X_16433_ CPU.registerFile\[12\]\[30\] _02826_ _02860_ _03901_ VGND VGND VPWR VPWR
+ _03902_ sky130_fd_sc_hd__o211a_1
X_10857_ net2356 _05708_ _06117_ VGND VGND VPWR VPWR _06126_ sky130_fd_sc_hd__mux2_1
X_13645_ CPU.registerFile\[15\]\[22\] _07236_ _07277_ CPU.registerFile\[11\]\[22\]
+ _07820_ VGND VGND VPWR VPWR _08066_ sky130_fd_sc_hd__o221a_1
XFILLER_0_156_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16364_ CPU.registerFile\[13\]\[28\] _02800_ VGND VGND VPWR VPWR _03835_ sky130_fd_sc_hd__or2_1
X_10788_ _06089_ VGND VGND VPWR VPWR _02108_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13576_ _07995_ _07998_ _07514_ VGND VGND VPWR VPWR _07999_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_143_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16593__64 clknet_1_0__leaf__03970_ VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__inv_2
X_18103_ net166 _02383_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15315_ _02813_ VGND VGND VPWR VPWR _02814_ sky130_fd_sc_hd__clkbuf_4
X_12527_ net2022 _04658_ _07085_ VGND VGND VPWR VPWR _07086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16295_ CPU.registerFile\[11\]\[26\] _02777_ VGND VGND VPWR VPWR _03768_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18034_ net1207 _02314_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_97_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12458_ _07048_ VGND VGND VPWR VPWR _07049_ sky130_fd_sc_hd__buf_4
XFILLER_0_140_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11409_ _05532_ net2050 _06419_ VGND VGND VPWR VPWR _06420_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12389_ _05488_ _06032_ VGND VGND VPWR VPWR _07012_ sky130_fd_sc_hd__nand2_2
XFILLER_0_50_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14128_ _08393_ VGND VGND VPWR VPWR _01472_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_128_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08620_ CPU.aluIn1\[19\] _04247_ VGND VGND VPWR VPWR _04340_ sky130_fd_sc_hd__or2_1
X_17818_ net1007 _02102_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_08551_ CPU.aluIn1\[8\] _04270_ VGND VGND VPWR VPWR _04271_ sky130_fd_sc_hd__or2_1
X_17749_ net938 _02033_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_141_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08482_ _04196_ _04197_ _04198_ VGND VGND VPWR VPWR _04202_ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09103_ _04782_ _04814_ net1277 VGND VGND VPWR VPWR _04815_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09034_ _04749_ VGND VGND VPWR VPWR _02577_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold320 per_uart.uart0.rx_count16\[0\] VGND VGND VPWR VPWR net1561 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold331 CPU.registerFile\[4\]\[29\] VGND VGND VPWR VPWR net1572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold342 CPU.registerFile\[6\]\[9\] VGND VGND VPWR VPWR net1583 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold353 CPU.registerFile\[6\]\[28\] VGND VGND VPWR VPWR net1594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 CPU.registerFile\[30\]\[25\] VGND VGND VPWR VPWR net1605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 CPU.registerFile\[16\]\[26\] VGND VGND VPWR VPWR net1616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold386 CPU.registerFile\[10\]\[30\] VGND VGND VPWR VPWR net1627 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold397 CPU.registerFile\[16\]\[4\] VGND VGND VPWR VPWR net1638 sky130_fd_sc_hd__dlygate4sd3_1
X_09936_ _05487_ net1620 _05559_ VGND VGND VPWR VPWR _05560_ sky130_fd_sc_hd__mux2_1
X_09867_ _05511_ net2394 _05512_ VGND VGND VPWR VPWR _05513_ sky130_fd_sc_hd__mux2_1
Xhold1020 CPU.registerFile\[27\]\[31\] VGND VGND VPWR VPWR net2261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1031 CPU.registerFile\[15\]\[31\] VGND VGND VPWR VPWR net2272 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1042 CPU.registerFile\[31\]\[2\] VGND VGND VPWR VPWR net2283 sky130_fd_sc_hd__dlygate4sd3_1
X_08818_ _04535_ _04536_ _04537_ VGND VGND VPWR VPWR _04538_ sky130_fd_sc_hd__a21o_1
Xhold1053 CPU.registerFile\[17\]\[21\] VGND VGND VPWR VPWR net2294 sky130_fd_sc_hd__dlygate4sd3_1
X_14508__630 clknet_1_1__leaf__02667_ VGND VGND VPWR VPWR net662 sky130_fd_sc_hd__inv_2
Xhold1064 CPU.registerFile\[24\]\[16\] VGND VGND VPWR VPWR net2305 sky130_fd_sc_hd__dlygate4sd3_1
X_09798_ net2355 _05109_ _05463_ VGND VGND VPWR VPWR _05470_ sky130_fd_sc_hd__mux2_1
Xhold1075 CPU.registerFile\[31\]\[21\] VGND VGND VPWR VPWR net2316 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1086 CPU.registerFile\[10\]\[14\] VGND VGND VPWR VPWR net2327 sky130_fd_sc_hd__dlygate4sd3_1
X_14965__1042 clknet_1_1__leaf__02712_ VGND VGND VPWR VPWR net1074 sky130_fd_sc_hd__inv_2
XANTENNA_204 _07841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1097 mapped_spi_flash.snd_bitcount\[5\] VGND VGND VPWR VPWR net2338 sky130_fd_sc_hd__dlygate4sd3_1
X_08749_ _04468_ _04233_ VGND VGND VPWR VPWR _04469_ sky130_fd_sc_hd__nor2_1
XANTENNA_215 _08302_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_226 clknet_1_1__leaf__02720_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_237 _02885_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_248 _03463_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11760_ _04714_ net2498 _06639_ VGND VGND VPWR VPWR _06642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_259 _05050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10711_ _05518_ net2000 _06045_ VGND VGND VPWR VPWR _06049_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11691_ net2490 _06590_ _06598_ _06594_ VGND VGND VPWR VPWR _01710_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13430_ CPU.registerFile\[31\]\[15\] _07347_ _07348_ CPU.registerFile\[27\]\[15\]
+ _07345_ VGND VGND VPWR VPWR _07858_ sky130_fd_sc_hd__o221a_1
X_10642_ _05843_ VGND VGND VPWR VPWR _06006_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13361_ _07519_ _07789_ _07790_ VGND VGND VPWR VPWR _07791_ sky130_fd_sc_hd__o21a_1
XFILLER_0_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10573_ net1320 mapped_spi_flash.rcv_bitcount\[4\] _05964_ VGND VGND VPWR VPWR _05965_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_64_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15100_ net1457 _07188_ VGND VGND VPWR VPWR _02737_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12312_ _06969_ VGND VGND VPWR VPWR _01426_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer9 net1251 VGND VGND VPWR VPWR net1250 sky130_fd_sc_hd__dlygate4sd1_1
X_16080_ CPU.registerFile\[26\]\[19\] _02861_ VGND VGND VPWR VPWR _03560_ sky130_fd_sc_hd__or2_1
X_13292_ CPU.registerFile\[31\]\[11\] _07403_ _07404_ CPU.registerFile\[27\]\[11\]
+ _07405_ VGND VGND VPWR VPWR _07724_ sky130_fd_sc_hd__o221a_1
XFILLER_0_122_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14554__672 clknet_1_1__leaf__02671_ VGND VGND VPWR VPWR net704 sky130_fd_sc_hd__inv_2
XFILLER_0_133_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12243_ CPU.aluIn1\[18\] _06916_ _06894_ VGND VGND VPWR VPWR _06917_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12174_ _06863_ _06864_ _06862_ VGND VGND VPWR VPWR _01493_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11125_ net2023 _05702_ _06263_ VGND VGND VPWR VPWR _06269_ sky130_fd_sc_hd__mux2_1
X_16982_ clknet_leaf_21_clk _01308_ VGND VGND VPWR VPWR CPU.rs2\[13\] sky130_fd_sc_hd__dfxtp_1
X_11056_ net2259 _05702_ _06226_ VGND VGND VPWR VPWR _06232_ sky130_fd_sc_hd__mux2_1
X_15933_ CPU.registerFile\[27\]\[15\] CPU.registerFile\[31\]\[15\] _02852_ VGND VGND
+ VPWR VPWR _03417_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10007_ net2004 _04696_ _05596_ VGND VGND VPWR VPWR _05598_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15864_ _03345_ _03349_ _03138_ VGND VGND VPWR VPWR _03350_ sky130_fd_sc_hd__a21o_1
X_17603_ net792 _01891_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_15795_ _03277_ _03282_ _03138_ VGND VGND VPWR VPWR _03283_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17534_ net723 _01822_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_106_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11958_ _05737_ _05489_ VGND VGND VPWR VPWR _06746_ sky130_fd_sc_hd__nand2_4
XFILLER_0_157_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10909_ _06142_ VGND VGND VPWR VPWR _06154_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17465_ net654 _01753_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[20\] sky130_fd_sc_hd__dfxtp_1
X_11889_ _06709_ VGND VGND VPWR VPWR _01624_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16416_ _03881_ _03885_ _02784_ VGND VGND VPWR VPWR _03886_ sky130_fd_sc_hd__a21o_1
XFILLER_0_156_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13628_ net1535 _08018_ _08049_ _08017_ VGND VGND VPWR VPWR _01316_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17396_ net585 _01684_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_14637__747 clknet_1_0__leaf__02679_ VGND VGND VPWR VPWR net779 sky130_fd_sc_hd__inv_2
XFILLER_0_54_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16347_ CPU.registerFile\[30\]\[27\] CPU.registerFile\[26\]\[27\] _03064_ VGND VGND
+ VPWR VPWR _03819_ sky130_fd_sc_hd__mux2_1
X_13559_ _07268_ _07979_ _07982_ VGND VGND VPWR VPWR _07983_ sky130_fd_sc_hd__or3_1
XFILLER_0_125_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16278_ _03750_ _03751_ _03317_ VGND VGND VPWR VPWR _03752_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18017_ net1190 _02297_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09721_ CPU.PC\[1\] _04872_ VGND VGND VPWR VPWR _05411_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_126_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14683__789 clknet_1_1__leaf__02683_ VGND VGND VPWR VPWR net821 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_143_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09652_ _05343_ _05344_ VGND VGND VPWR VPWR _05345_ sky130_fd_sc_hd__xor2_1
X_14382__517 clknet_1_1__leaf__02654_ VGND VGND VPWR VPWR net549 sky130_fd_sc_hd__inv_2
X_08603_ _04321_ _04322_ VGND VGND VPWR VPWR _04323_ sky130_fd_sc_hd__nor2_1
XFILLER_0_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09583_ mapped_spi_ram.rcv_data\[30\] net17 _04643_ per_uart.rx_data\[6\] VGND VGND
+ VPWR VPWR _05278_ sky130_fd_sc_hd__a22o_1
X_08534_ CPU.rs2\[16\] _04200_ _04205_ VGND VGND VPWR VPWR _04254_ sky130_fd_sc_hd__a21o_2
XFILLER_0_77_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16557__31 clknet_1_1__leaf__03967_ VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__inv_2
XFILLER_0_46_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16572__45 clknet_1_1__leaf__03968_ VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_21_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_154_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09017_ _04463_ _04465_ _04353_ VGND VGND VPWR VPWR _04733_ sky130_fd_sc_hd__a21oi_1
Xhold150 mapped_spi_flash.cmd_addr\[8\] VGND VGND VPWR VPWR net1391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 mapped_spi_flash.cmd_addr\[4\] VGND VGND VPWR VPWR net1402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 _01722_ VGND VGND VPWR VPWR net1413 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold183 mapped_spi_ram.rcv_data\[16\] VGND VGND VPWR VPWR net1424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold194 mapped_spi_ram.rcv_data\[17\] VGND VGND VPWR VPWR net1435 sky130_fd_sc_hd__dlygate4sd3_1
X_09919_ _05547_ net2451 _05533_ VGND VGND VPWR VPWR _05548_ sky130_fd_sc_hd__mux2_1
X_12930_ _07370_ VGND VGND VPWR VPWR _07371_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ mapped_spi_ram.rcv_data\[15\] _04689_ _04691_ mapped_spi_flash.rcv_data\[15\]
+ VGND VGND VPWR VPWR _07304_ sky130_fd_sc_hd__a22o_2
XFILLER_0_158_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11812_ _05359_ net2120 _06661_ VGND VGND VPWR VPWR _06669_ sky130_fd_sc_hd__mux2_1
X_15580_ _05439_ VGND VGND VPWR VPWR _03074_ sky130_fd_sc_hd__clkbuf_4
X_12792_ _07234_ VGND VGND VPWR VPWR _07235_ sky130_fd_sc_hd__buf_2
XFILLER_0_84_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11743_ net1344 _06570_ VGND VGND VPWR VPWR _06631_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17250_ net440 _01538_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14462_ clknet_1_1__leaf__02653_ VGND VGND VPWR VPWR _02662_ sky130_fd_sc_hd__buf_1
X_11674_ mapped_spi_ram.rcv_data\[22\] _06588_ VGND VGND VPWR VPWR _06589_ sky130_fd_sc_hd__or2_1
X_15169__1195 clknet_1_1__leaf__02747_ VGND VGND VPWR VPWR net1227 sky130_fd_sc_hd__inv_2
X_16201_ _02898_ _03674_ _03675_ _03676_ _02887_ VGND VGND VPWR VPWR _03677_ sky130_fd_sc_hd__o221a_1
XFILLER_0_138_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13413_ _07837_ _07840_ _07320_ VGND VGND VPWR VPWR _07841_ sky130_fd_sc_hd__mux2_2
XFILLER_0_154_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17181_ clknet_leaf_24_clk _01469_ VGND VGND VPWR VPWR CPU.Bimm\[4\] sky130_fd_sc_hd__dfxtp_1
X_10625_ mapped_spi_flash.rcv_data\[11\] _05994_ VGND VGND VPWR VPWR _05997_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16132_ CPU.registerFile\[24\]\[21\] _03130_ _02780_ _03609_ VGND VGND VPWR VPWR
+ _03610_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_77_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13344_ CPU.registerFile\[8\]\[13\] CPU.registerFile\[12\]\[13\] _07233_ VGND VGND
+ VPWR VPWR _07774_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10556_ mapped_spi_flash.snd_bitcount\[4\] _05944_ VGND VGND VPWR VPWR _05953_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16063_ _02901_ _03541_ _03542_ _03030_ VGND VGND VPWR VPWR _03543_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10487_ net1383 _05887_ _05851_ _05896_ VGND VGND VPWR VPWR _05897_ sky130_fd_sc_hd__a211o_1
X_13275_ _07364_ _07706_ VGND VGND VPWR VPWR _07707_ sky130_fd_sc_hd__or2_1
X_12226_ CPU.aluIn1\[22\] _06903_ _06894_ VGND VGND VPWR VPWR _06904_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14218__394 clknet_1_1__leaf__08431_ VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__inv_2
X_12157_ _06851_ VGND VGND VPWR VPWR _01497_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_9_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11108_ net2360 _05685_ _06252_ VGND VGND VPWR VPWR _06260_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16965_ net260 _01291_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_12088_ _05402_ net2008 _06805_ VGND VGND VPWR VPWR _06815_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_108_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15916_ CPU.registerFile\[8\]\[15\] CPU.registerFile\[12\]\[15\] _02798_ VGND VGND
+ VPWR VPWR _03400_ sky130_fd_sc_hd__mux2_1
X_11039_ net1882 _05685_ _06215_ VGND VGND VPWR VPWR _06223_ sky130_fd_sc_hd__mux2_1
X_16896_ _04644_ _06468_ VGND VGND VPWR VPWR _04174_ sky130_fd_sc_hd__nand2_1
X_15847_ CPU.registerFile\[14\]\[13\] CPU.registerFile\[10\]\[13\] _03082_ VGND VGND
+ VPWR VPWR _03333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_121_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15778_ CPU.registerFile\[12\]\[11\] _03118_ VGND VGND VPWR VPWR _03266_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17517_ net706 _01805_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_14729_ clknet_1_0__leaf__02686_ VGND VGND VPWR VPWR _02689_ sky130_fd_sc_hd__buf_1
XFILLER_0_47_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17448_ net637 _01736_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17379_ net568 _01667_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_136_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14964__1041 clknet_1_1__leaf__02712_ VGND VGND VPWR VPWR net1073 sky130_fd_sc_hd__inv_2
XFILLER_0_2_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_151_Right_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09704_ net1294 _05394_ VGND VGND VPWR VPWR _05395_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_52_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09635_ _05328_ _04880_ VGND VGND VPWR VPWR _05329_ sky130_fd_sc_hd__xnor2_1
X_09566_ _04278_ _04312_ _04275_ VGND VGND VPWR VPWR _05262_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08517_ CPU.rs2\[23\] _04201_ _04206_ VGND VGND VPWR VPWR _04237_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09497_ CPU.PC\[9\] _04920_ CPU.PC\[10\] VGND VGND VPWR VPWR _05196_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_156_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10410_ _05836_ VGND VGND VPWR VPWR _02232_ sky130_fd_sc_hd__clkbuf_1
X_11390_ _05514_ net1771 _06408_ VGND VGND VPWR VPWR _06410_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_59_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10341_ _05518_ net2244 _05788_ VGND VGND VPWR VPWR _05792_ sky130_fd_sc_hd__mux2_1
X_13060_ CPU.registerFile\[18\]\[5\] CPU.registerFile\[22\]\[5\] _07314_ VGND VGND
+ VPWR VPWR _07498_ sky130_fd_sc_hd__mux2_1
X_10272_ _05518_ net1741 _05751_ VGND VGND VPWR VPWR _05755_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12011_ _06774_ VGND VGND VPWR VPWR _01567_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_72_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14666__773 clknet_1_1__leaf__02682_ VGND VGND VPWR VPWR net805 sky130_fd_sc_hd__inv_2
X_16750_ _05096_ _08454_ _05288_ VGND VGND VPWR VPWR _04068_ sky130_fd_sc_hd__and3b_1
X_15701_ net2496 _03081_ _03191_ _03080_ VGND VGND VPWR VPWR _02422_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12913_ _07344_ _07346_ _07350_ _07354_ _07302_ VGND VGND VPWR VPWR _07355_ sky130_fd_sc_hd__a221o_1
X_16681_ _04004_ _04009_ _06030_ VGND VGND VPWR VPWR _02584_ sky130_fd_sc_hd__a21oi_1
X_13893_ CPU.registerFile\[5\]\[30\] CPU.registerFile\[4\]\[30\] _04985_ VGND VGND
+ VPWR VPWR _08306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15632_ CPU.registerFile\[13\]\[7\] _03123_ VGND VGND VPWR VPWR _03124_ sky130_fd_sc_hd__or2_1
X_12844_ CPU.registerFile\[13\]\[0\] _07282_ _07286_ VGND VGND VPWR VPWR _07287_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_103_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18351_ clknet_leaf_1_clk _02631_ VGND VGND VPWR VPWR per_uart.uart0.rx_bitcount\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_15563_ _08395_ VGND VGND VPWR VPWR _03057_ sky130_fd_sc_hd__buf_4
XFILLER_0_57_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14064__339 clknet_1_1__leaf__08366_ VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__inv_2
XFILLER_0_56_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17302_ net491 _01590_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11726_ net1308 mapped_spi_ram.div_counter\[1\] VGND VGND VPWR VPWR _06618_ sky130_fd_sc_hd__nand2_1
X_18282_ net115 _02562_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_15494_ CPU.registerFile\[18\]\[3\] _02832_ _02835_ CPU.registerFile\[19\]\[3\] _02796_
+ VGND VGND VPWR VPWR _02990_ sky130_fd_sc_hd__o221a_1
XFILLER_0_84_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_801 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_140_Left_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17233_ net423 _01521_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_16536__12 clknet_1_1__leaf__03965_ VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__inv_2
Xclkbuf_0__03971_ _03971_ VGND VGND VPWR VPWR clknet_0__03971_ sky130_fd_sc_hd__clkbuf_16
X_11657_ net1407 _06575_ _06579_ _06539_ VGND VGND VPWR VPWR _01725_ sky130_fd_sc_hd__o211a_1
X_14831__921 clknet_1_1__leaf__02699_ VGND VGND VPWR VPWR net953 sky130_fd_sc_hd__inv_2
XFILLER_0_126_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17164_ net388 _01452_ VGND VGND VPWR VPWR CPU.aluReg\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10608_ net1458 _05981_ VGND VGND VPWR VPWR _05987_ sky130_fd_sc_hd__or2_1
X_11588_ net1406 _06524_ _06530_ _06516_ VGND VGND VPWR VPWR _01745_ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16115_ CPU.registerFile\[26\]\[20\] _02861_ VGND VGND VPWR VPWR _03594_ sky130_fd_sc_hd__or2_1
X_13327_ _07519_ _07756_ _07757_ VGND VGND VPWR VPWR _07758_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold908 CPU.registerFile\[6\]\[16\] VGND VGND VPWR VPWR net2149 sky130_fd_sc_hd__dlygate4sd3_1
X_16551__26 clknet_1_1__leaf__03966_ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__inv_2
X_17095_ net353 _01417_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[25\] sky130_fd_sc_hd__dfxtp_1
Xhold919 CPU.registerFile\[29\]\[31\] VGND VGND VPWR VPWR net2160 sky130_fd_sc_hd__dlygate4sd3_1
X_10539_ mapped_spi_flash.cmd_addr\[0\] _05824_ _05827_ mapped_spi_flash.cmd_addr\[1\]
+ VGND VGND VPWR VPWR _05939_ sky130_fd_sc_hd__a22o_1
Xclkbuf_1_1__f__02753_ clknet_0__02753_ VGND VGND VPWR VPWR clknet_1_1__leaf__02753_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0__08360_ _08360_ VGND VGND VPWR VPWR clknet_0__08360_ sky130_fd_sc_hd__clkbuf_16
X_16046_ _02926_ _03525_ _03526_ VGND VGND VPWR VPWR _03527_ sky130_fd_sc_hd__o21a_1
X_13258_ _07412_ _07689_ _07690_ VGND VGND VPWR VPWR _07691_ sky130_fd_sc_hd__o21a_1
X_14749__848 clknet_1_1__leaf__02690_ VGND VGND VPWR VPWR net880 sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__02684_ clknet_0__02684_ VGND VGND VPWR VPWR clknet_1_1__leaf__02684_
+ sky130_fd_sc_hd__clkbuf_16
X_12209_ _06861_ VGND VGND VPWR VPWR _06891_ sky130_fd_sc_hd__clkbuf_4
X_13189_ CPU.registerFile\[8\]\[8\] CPU.registerFile\[12\]\[8\] _07315_ VGND VGND
+ VPWR VPWR _07624_ sky130_fd_sc_hd__mux2_1
X_16509__178 clknet_1_0__leaf__03962_ VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__inv_2
X_17997_ clknet_leaf_8_clk _02281_ VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[11\]
+ sky130_fd_sc_hd__dfxtp_1
X_16948_ net243 _01274_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_16879_ _04193_ _04158_ _04161_ _04162_ VGND VGND VPWR VPWR _04163_ sky130_fd_sc_hd__and4_1
X_09420_ _05117_ _05122_ _04773_ VGND VGND VPWR VPWR _05123_ sky130_fd_sc_hd__o21a_1
X_09351_ _04800_ _05054_ _05056_ _04678_ VGND VGND VPWR VPWR _05057_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09282_ _04341_ _04683_ VGND VGND VPWR VPWR _04991_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_23_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14494__618 clknet_1_1__leaf__02665_ VGND VGND VPWR VPWR net650 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_138_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_151_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload70 clknet_1_1__leaf__02677_ VGND VGND VPWR VPWR clkload70/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_3_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14234__409 clknet_1_1__leaf__08432_ VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__inv_2
Xclkload81 clknet_1_1__leaf__02663_ VGND VGND VPWR VPWR clkload81/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_140_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload92 clknet_1_0__leaf__08467_ VGND VGND VPWR VPWR clkload92/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_11_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14808__901 clknet_1_1__leaf__02696_ VGND VGND VPWR VPWR net933 sky130_fd_sc_hd__inv_2
XFILLER_0_100_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08997_ net1665 _04714_ _04668_ VGND VGND VPWR VPWR _04715_ sky130_fd_sc_hd__mux2_1
X_15168__1194 clknet_1_0__leaf__02747_ VGND VGND VPWR VPWR net1226 sky130_fd_sc_hd__inv_2
X_12748__201 clknet_1_0__leaf__07221_ VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_149_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09618_ _05308_ _05280_ _05310_ _05311_ _04716_ VGND VGND VPWR VPWR _05312_ sky130_fd_sc_hd__a221o_1
X_15215__126 clknet_1_0__leaf__02752_ VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__inv_2
X_10890_ _06144_ VGND VGND VPWR VPWR _02061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09549_ _04426_ _04404_ _04425_ VGND VGND VPWR VPWR _05246_ sky130_fd_sc_hd__nor3_1
XFILLER_0_65_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12560_ net2519 _05108_ _07096_ VGND VGND VPWR VPWR _07103_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_778 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11511_ net1398 _06473_ _06476_ VGND VGND VPWR VPWR _06477_ sky130_fd_sc_hd__a21oi_1
X_12491_ _07066_ VGND VGND VPWR VPWR _01344_ sky130_fd_sc_hd__clkbuf_1
X_11442_ _06437_ VGND VGND VPWR VPWR _01802_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14161_ _08417_ VGND VGND VPWR VPWR _01481_ sky130_fd_sc_hd__clkbuf_1
X_11373_ _05497_ CPU.registerFile\[24\]\[28\] _06397_ VGND VGND VPWR VPWR _06401_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13112_ CPU.registerFile\[9\]\[6\] _07503_ _07548_ _07296_ _07349_ VGND VGND VPWR
+ VPWR _07549_ sky130_fd_sc_hd__o221a_1
X_10324_ _05501_ net2062 _05777_ VGND VGND VPWR VPWR _05783_ sky130_fd_sc_hd__mux2_1
X_14092_ _05311_ _08369_ _08371_ _08372_ VGND VGND VPWR VPWR _08373_ sky130_fd_sc_hd__and4_1
XFILLER_0_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13043_ _07235_ VGND VGND VPWR VPWR _07482_ sky130_fd_sc_hd__buf_4
X_10255_ _05501_ net2473 _05740_ VGND VGND VPWR VPWR _05746_ sky130_fd_sc_hd__mux2_1
X_17920_ net1109 _02204_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[0\] sky130_fd_sc_hd__dfxtp_1
X_17851_ net1040 _02135_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_10186_ _05065_ VGND VGND VPWR VPWR _05700_ sky130_fd_sc_hd__clkbuf_4
X_16802_ net5 net1536 _04193_ VGND VGND VPWR VPWR _04111_ sky130_fd_sc_hd__mux2_1
X_17782_ net971 _02066_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_16733_ _03995_ _05158_ _07132_ VGND VGND VPWR VPWR _04054_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13945_ net1341 _08355_ _05855_ VGND VGND VPWR VPWR _01327_ sky130_fd_sc_hd__o21ai_1
X_16664_ _05289_ VGND VGND VPWR VPWR _03995_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_85_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13876_ CPU.registerFile\[28\]\[29\] CPU.registerFile\[24\]\[29\] _07297_ VGND VGND
+ VPWR VPWR _08290_ sky130_fd_sc_hd__mux2_1
X_14963__1040 clknet_1_1__leaf__02712_ VGND VGND VPWR VPWR net1072 sky130_fd_sc_hd__inv_2
XFILLER_0_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15615_ CPU.registerFile\[18\]\[6\] _02833_ _02836_ CPU.registerFile\[19\]\[6\] _02758_
+ VGND VGND VPWR VPWR _03108_ sky130_fd_sc_hd__o221a_1
XFILLER_0_9_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12827_ _07232_ _07251_ _07269_ VGND VGND VPWR VPWR _07270_ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18334_ clknet_leaf_7_clk _02614_ VGND VGND VPWR VPWR per_uart.uart0.tx_bitcount\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_15546_ _02759_ _03037_ _03039_ _02767_ VGND VGND VPWR VPWR _03040_ sky130_fd_sc_hd__a211o_1
X_12758_ clknet_1_1__leaf__07222_ VGND VGND VPWR VPWR _07223_ sky130_fd_sc_hd__buf_1
XFILLER_0_45_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11709_ mapped_spi_ram.rcv_data\[7\] _06601_ VGND VGND VPWR VPWR _06609_ sky130_fd_sc_hd__or2_1
X_18265_ clknet_leaf_2_clk _02545_ VGND VGND VPWR VPWR per_uart.uart0.rxd_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_15477_ CPU.registerFile\[29\]\[3\] _02926_ VGND VGND VPWR VPWR _02973_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12689_ _07172_ net1422 VGND VGND VPWR VPWR _00036_ sky130_fd_sc_hd__nor2_1
X_17216_ net406 _01504_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18196_ net227 _02476_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17147_ net371 _01435_ VGND VGND VPWR VPWR CPU.aluReg\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_116_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold705 CPU.registerFile\[25\]\[20\] VGND VGND VPWR VPWR net1946 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold716 CPU.registerFile\[26\]\[9\] VGND VGND VPWR VPWR net1957 sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 CPU.registerFile\[22\]\[22\] VGND VGND VPWR VPWR net1968 sky130_fd_sc_hd__dlygate4sd3_1
X_14337__477 clknet_1_1__leaf__08466_ VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__inv_2
Xhold738 CPU.registerFile\[7\]\[2\] VGND VGND VPWR VPWR net1979 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17078_ net336 _01400_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[8\] sky130_fd_sc_hd__dfxtp_1
Xhold749 CPU.registerFile\[19\]\[11\] VGND VGND VPWR VPWR net1990 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16029_ _02911_ _03507_ _03509_ _03245_ VGND VGND VPWR VPWR _03510_ sky130_fd_sc_hd__a211o_1
X_08920_ CPU.PC\[1\] _04598_ _04637_ _04590_ _04639_ VGND VGND VPWR VPWR _04640_ sky130_fd_sc_hd__a221oi_1
X_13975__259 clknet_1_1__leaf__08357_ VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__02667_ clknet_0__02667_ VGND VGND VPWR VPWR clknet_1_1__leaf__02667_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08851_ _04568_ _04565_ _04564_ _04569_ _04570_ VGND VGND VPWR VPWR _04571_ sky130_fd_sc_hd__o311a_4
Xclkbuf_0__02698_ _02698_ VGND VGND VPWR VPWR clknet_0__02698_ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_0__07225_ _07225_ VGND VGND VPWR VPWR clknet_0__07225_ sky130_fd_sc_hd__clkbuf_16
X_08782_ _04501_ VGND VGND VPWR VPWR _04502_ sky130_fd_sc_hd__buf_1
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14803__897 clknet_1_0__leaf__02695_ VGND VGND VPWR VPWR net929 sky130_fd_sc_hd__inv_2
XFILLER_0_67_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09403_ _05103_ _05104_ _05106_ _04492_ VGND VGND VPWR VPWR _05107_ sky130_fd_sc_hd__o31a_2
XFILLER_0_48_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14047__323 clknet_1_1__leaf__08365_ VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__inv_2
X_14502__625 clknet_1_1__leaf__02666_ VGND VGND VPWR VPWR net657 sky130_fd_sc_hd__inv_2
X_09334_ _04837_ _04903_ VGND VGND VPWR VPWR _05041_ sky130_fd_sc_hd__and2b_1
X_14240__413 clknet_1_0__leaf__08434_ VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__inv_2
XFILLER_0_63_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12778__227 clknet_1_1__leaf__07225_ VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__inv_2
X_09265_ _04825_ _04907_ VGND VGND VPWR VPWR _04975_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09196_ _04825_ _04907_ _04823_ VGND VGND VPWR VPWR _04908_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10040_ net2256 _05130_ _05607_ VGND VGND VPWR VPWR _05615_ sky130_fd_sc_hd__mux2_1
Xhold76 _02197_ VGND VGND VPWR VPWR net1317 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 CPU.cycles\[0\] VGND VGND VPWR VPWR net1328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 per_uart.uart0.enable16_counter\[3\] VGND VGND VPWR VPWR net1339 sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ _05090_ net2077 _06758_ VGND VGND VPWR VPWR _06764_ sky130_fd_sc_hd__mux2_1
X_13730_ CPU.registerFile\[25\]\[25\] CPU.registerFile\[29\]\[25\] _05284_ VGND VGND
+ VPWR VPWR _08148_ sky130_fd_sc_hd__mux2_1
X_10942_ _06171_ VGND VGND VPWR VPWR _02036_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_67_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__02756_ clknet_0__02756_ VGND VGND VPWR VPWR clknet_1_0__leaf__02756_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14778__874 clknet_1_0__leaf__02693_ VGND VGND VPWR VPWR net906 sky130_fd_sc_hd__inv_2
X_13661_ CPU.registerFile\[26\]\[23\] _07801_ _04987_ _08080_ VGND VGND VPWR VPWR
+ _08081_ sky130_fd_sc_hd__o211a_1
X_10873_ _06134_ VGND VGND VPWR VPWR _02068_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__02687_ clknet_0__02687_ VGND VGND VPWR VPWR clknet_1_0__leaf__02687_
+ sky130_fd_sc_hd__clkbuf_16
X_15400_ _04620_ VGND VGND VPWR VPWR _02898_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_155_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12612_ _07122_ _07128_ _07129_ _07121_ VGND VGND VPWR VPWR _00003_ sky130_fd_sc_hd__o22ai_1
X_16380_ CPU.registerFile\[2\]\[28\] _02821_ _02813_ CPU.registerFile\[3\]\[28\] _05070_
+ VGND VGND VPWR VPWR _03851_ sky130_fd_sc_hd__a221o_1
X_13592_ _07308_ VGND VGND VPWR VPWR _08015_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_155_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15331_ CPU.registerFile\[22\]\[0\] CPU.registerFile\[23\]\[0\] _02829_ VGND VGND
+ VPWR VPWR _02830_ sky130_fd_sc_hd__mux2_1
X_12543_ net2528 _04932_ _07085_ VGND VGND VPWR VPWR _07094_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18050_ net1223 _02330_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15262_ _02760_ VGND VGND VPWR VPWR _02761_ sky130_fd_sc_hd__clkbuf_8
X_12474_ _07057_ VGND VGND VPWR VPWR _01352_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17001_ clknet_leaf_11_clk _00001_ VGND VGND VPWR VPWR CPU.state\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14213_ clknet_1_0__leaf__08363_ VGND VGND VPWR VPWR _08431_ sky130_fd_sc_hd__buf_1
XFILLER_0_123_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11425_ _05549_ CPU.registerFile\[24\]\[3\] _06419_ VGND VGND VPWR VPWR _06428_ sky130_fd_sc_hd__mux2_1
XANTENNA_7 _02807_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14144_ _08406_ VGND VGND VPWR VPWR _01475_ sky130_fd_sc_hd__clkbuf_1
X_11356_ _05549_ net2390 _06382_ VGND VGND VPWR VPWR _06391_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10307_ _05553_ net2027 _05739_ VGND VGND VPWR VPWR _05773_ sky130_fd_sc_hd__mux2_1
X_11287_ _06354_ VGND VGND VPWR VPWR _01874_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_111_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13026_ _07360_ _07460_ _07464_ _07380_ VGND VGND VPWR VPWR _07465_ sky130_fd_sc_hd__o211a_1
X_17903_ net1092 net1325 VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[21\] sky130_fd_sc_hd__dfxtp_1
X_10238_ _05447_ VGND VGND VPWR VPWR _05735_ sky130_fd_sc_hd__clkbuf_4
X_10169_ _05688_ VGND VGND VPWR VPWR _02341_ sky130_fd_sc_hd__clkbuf_1
X_17834_ net1023 _02118_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_17765_ net954 _02049_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer19 net1261 VGND VGND VPWR VPWR net1260 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_16_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13928_ CPU.registerFile\[14\]\[31\] CPU.registerFile\[10\]\[31\] _07480_ VGND VGND
+ VPWR VPWR _08340_ sky130_fd_sc_hd__mux2_1
X_16716_ _08453_ VGND VGND VPWR VPWR _04039_ sky130_fd_sc_hd__buf_2
XFILLER_0_89_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17696_ net885 _01984_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13859_ CPU.registerFile\[18\]\[29\] CPU.registerFile\[22\]\[29\] _07785_ VGND VGND
+ VPWR VPWR _08273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_851 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18317_ clknet_leaf_16_clk _02597_ VGND VGND VPWR VPWR CPU.PC\[17\] sky130_fd_sc_hd__dfxtp_1
X_15529_ CPU.registerFile\[22\]\[4\] _08399_ VGND VGND VPWR VPWR _03024_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_33_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09050_ _04353_ _04463_ _04465_ VGND VGND VPWR VPWR _04764_ sky130_fd_sc_hd__and3_1
X_15167__1193 clknet_1_0__leaf__02747_ VGND VGND VPWR VPWR net1225 sky130_fd_sc_hd__inv_2
X_18248_ net89 _02528_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18179_ net210 _02459_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold502 CPU.registerFile\[19\]\[30\] VGND VGND VPWR VPWR net1743 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold513 CPU.registerFile\[27\]\[25\] VGND VGND VPWR VPWR net1754 sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 CPU.registerFile\[6\]\[18\] VGND VGND VPWR VPWR net1765 sky130_fd_sc_hd__dlygate4sd3_1
X_15244__152 clknet_1_1__leaf__02755_ VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__inv_2
XFILLER_0_12_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold535 CPU.registerFile\[17\]\[20\] VGND VGND VPWR VPWR net1776 sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 CPU.registerFile\[2\]\[27\] VGND VGND VPWR VPWR net1787 sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 _04146_ VGND VGND VPWR VPWR net1798 sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 CPU.registerFile\[19\]\[23\] VGND VGND VPWR VPWR net1809 sky130_fd_sc_hd__dlygate4sd3_1
X_09952_ _05507_ net1629 _05559_ VGND VGND VPWR VPWR _05568_ sky130_fd_sc_hd__mux2_1
Xhold579 CPU.PC\[11\] VGND VGND VPWR VPWR net1820 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08903_ CPU.aluIn1\[0\] _04523_ VGND VGND VPWR VPWR _04623_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09883_ _05523_ VGND VGND VPWR VPWR _02494_ sky130_fd_sc_hd__clkbuf_1
Xhold1202 CPU.registerFile\[8\]\[25\] VGND VGND VPWR VPWR net2443 sky130_fd_sc_hd__dlygate4sd3_1
X_08834_ CPU.aluIn1\[15\] _04494_ VGND VGND VPWR VPWR _04554_ sky130_fd_sc_hd__xnor2_2
Xhold1213 CPU.registerFile\[23\]\[6\] VGND VGND VPWR VPWR net2454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1224 CPU.registerFile\[24\]\[7\] VGND VGND VPWR VPWR net2465 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1235 CPU.aluIn1\[31\] VGND VGND VPWR VPWR net2476 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1246 CPU.registerFile\[14\]\[5\] VGND VGND VPWR VPWR net2487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1257 CPU.registerFile\[13\]\[29\] VGND VGND VPWR VPWR net2498 sky130_fd_sc_hd__dlygate4sd3_1
X_08765_ _04483_ _04484_ VGND VGND VPWR VPWR _04485_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1268 mapped_spi_ram.rcv_data\[12\] VGND VGND VPWR VPWR net2509 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1279 CPU.registerFile\[13\]\[27\] VGND VGND VPWR VPWR net2520 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_408 _04659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_419 _03296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08696_ _04410_ _04414_ _04415_ VGND VGND VPWR VPWR _04416_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_49_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09317_ _04818_ _05022_ _05024_ _04916_ VGND VGND VPWR VPWR _05025_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_62_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09248_ net2147 _04958_ _04668_ VGND VGND VPWR VPWR _04959_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09179_ _04857_ _04889_ _04890_ VGND VGND VPWR VPWR _04891_ sky130_fd_sc_hd__o21a_1
XFILLER_0_121_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11210_ _05539_ net1961 _06310_ VGND VGND VPWR VPWR _06314_ sky130_fd_sc_hd__mux2_1
X_12190_ _06876_ VGND VGND VPWR VPWR _01455_ sky130_fd_sc_hd__clkbuf_1
Xoutput11 net11 VGND VGND VPWR VPWR spi_mosi sky130_fd_sc_hd__buf_2
Xoutput9 net9 VGND VGND VPWR VPWR spi_cs_n sky130_fd_sc_hd__buf_2
X_11141_ _06277_ VGND VGND VPWR VPWR _01943_ sky130_fd_sc_hd__clkbuf_1
X_13958__243 clknet_1_0__leaf__08356_ VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__inv_2
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11072_ _06240_ VGND VGND VPWR VPWR _01975_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14019__299 clknet_1_0__leaf__08361_ VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__inv_2
X_10023_ net2101 _04958_ _05596_ VGND VGND VPWR VPWR _05606_ sky130_fd_sc_hd__mux2_1
X_15880_ CPU.aluIn1\[13\] _03081_ _03365_ _03080_ VGND VGND VPWR VPWR _02427_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14212__389 clknet_1_1__leaf__08430_ VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__inv_2
XFILLER_0_53_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17550_ net739 _01838_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_14762_ clknet_1_1__leaf__02686_ VGND VGND VPWR VPWR _02692_ sky130_fd_sc_hd__buf_1
X_11974_ _04798_ net2002 _06747_ VGND VGND VPWR VPWR _06755_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13713_ CPU.registerFile\[9\]\[24\] _07383_ _08131_ VGND VGND VPWR VPWR _08132_ sky130_fd_sc_hd__o21a_1
X_10925_ _06162_ VGND VGND VPWR VPWR _02044_ sky130_fd_sc_hd__clkbuf_1
X_17481_ net670 net27 VGND VGND VPWR VPWR mapped_spi_flash.div_counter\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16432_ CPU.registerFile\[8\]\[30\] _02777_ VGND VGND VPWR VPWR _03901_ sky130_fd_sc_hd__or2_1
XFILLER_0_156_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13644_ CPU.registerFile\[14\]\[22\] CPU.registerFile\[10\]\[22\] _07480_ VGND VGND
+ VPWR VPWR _08065_ sky130_fd_sc_hd__mux2_1
X_10856_ _06125_ VGND VGND VPWR VPWR _02076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16363_ CPU.registerFile\[15\]\[28\] CPU.registerFile\[11\]\[28\] _02906_ VGND VGND
+ VPWR VPWR _03834_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13575_ _07650_ _07996_ _07997_ VGND VGND VPWR VPWR _07998_ sky130_fd_sc_hd__o21ai_2
X_10787_ _05526_ net1896 _06081_ VGND VGND VPWR VPWR _06089_ sky130_fd_sc_hd__mux2_1
X_18102_ net165 _02382_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_30_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15314_ net15 _05405_ VGND VGND VPWR VPWR _02813_ sky130_fd_sc_hd__nor2_2
X_12526_ _07084_ VGND VGND VPWR VPWR _07085_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_81_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16294_ CPU.registerFile\[9\]\[26\] CPU.registerFile\[13\]\[26\] _02999_ VGND VGND
+ VPWR VPWR _03767_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18033_ net1206 _02313_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[27\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_97_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12457_ _05450_ _05669_ VGND VGND VPWR VPWR _07048_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_113_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11408_ _06396_ VGND VGND VPWR VPWR _06419_ sky130_fd_sc_hd__clkbuf_4
X_12388_ _07011_ VGND VGND VPWR VPWR _01392_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14127_ _04483_ _05111_ _08387_ VGND VGND VPWR VPWR _08393_ sky130_fd_sc_hd__mux2_1
X_14531__651 clknet_1_1__leaf__02669_ VGND VGND VPWR VPWR net683 sky130_fd_sc_hd__inv_2
X_11339_ _06359_ VGND VGND VPWR VPWR _06382_ sky130_fd_sc_hd__buf_4
XFILLER_0_120_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13009_ _07291_ _07448_ VGND VGND VPWR VPWR _07449_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_128_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14449__578 clknet_1_0__leaf__02660_ VGND VGND VPWR VPWR net610 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_128_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17817_ net1006 _02101_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_08550_ CPU.rs2\[8\] CPU.Bimm\[8\] net1295 VGND VGND VPWR VPWR _04270_ sky130_fd_sc_hd__mux2_1
X_14187__366 clknet_1_0__leaf__08428_ VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__inv_2
X_17748_ net937 _02032_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08481_ _04200_ VGND VGND VPWR VPWR _04201_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_141_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17679_ net868 _01967_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09102_ _04648_ VGND VGND VPWR VPWR _04814_ sky130_fd_sc_hd__buf_4
XFILLER_0_150_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14915__998 clknet_1_0__leaf__02706_ VGND VGND VPWR VPWR net1030 sky130_fd_sc_hd__inv_2
XFILLER_0_127_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09033_ net1613 _04748_ _04668_ VGND VGND VPWR VPWR _04749_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14614__726 clknet_1_1__leaf__02677_ VGND VGND VPWR VPWR net758 sky130_fd_sc_hd__inv_2
XFILLER_0_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold310 mapped_spi_flash.clk_div VGND VGND VPWR VPWR net1551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 CPU.PC\[3\] VGND VGND VPWR VPWR net1562 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold332 CPU.registerFile\[5\]\[17\] VGND VGND VPWR VPWR net1573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold343 CPU.registerFile\[5\]\[3\] VGND VGND VPWR VPWR net1584 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold354 CPU.registerFile\[5\]\[13\] VGND VGND VPWR VPWR net1595 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold365 CPU.registerFile\[9\]\[25\] VGND VGND VPWR VPWR net1606 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 CPU.registerFile\[7\]\[27\] VGND VGND VPWR VPWR net1617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 CPU.registerFile\[9\]\[26\] VGND VGND VPWR VPWR net1628 sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 CPU.registerFile\[2\]\[30\] VGND VGND VPWR VPWR net1639 sky130_fd_sc_hd__dlygate4sd3_1
X_09935_ _05558_ VGND VGND VPWR VPWR _05559_ sky130_fd_sc_hd__buf_4
X_09866_ _05490_ VGND VGND VPWR VPWR _05512_ sky130_fd_sc_hd__buf_4
Xhold1010 CPU.registerFile\[10\]\[21\] VGND VGND VPWR VPWR net2251 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 per_uart.d_in_uart\[6\] VGND VGND VPWR VPWR net2262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1032 CPU.registerFile\[10\]\[25\] VGND VGND VPWR VPWR net2273 sky130_fd_sc_hd__dlygate4sd3_1
X_08817_ CPU.aluIn1\[5\] CPU.Bimm\[5\] VGND VGND VPWR VPWR _04537_ sky130_fd_sc_hd__and2_1
Xhold1043 CPU.registerFile\[12\]\[29\] VGND VGND VPWR VPWR net2284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1054 CPU.registerFile\[22\]\[27\] VGND VGND VPWR VPWR net2295 sky130_fd_sc_hd__dlygate4sd3_1
X_09797_ _05469_ VGND VGND VPWR VPWR _02526_ sky130_fd_sc_hd__clkbuf_1
Xhold1065 CPU.registerFile\[18\]\[10\] VGND VGND VPWR VPWR net2306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1076 CPU.registerFile\[18\]\[27\] VGND VGND VPWR VPWR net2317 sky130_fd_sc_hd__dlygate4sd3_1
X_08748_ CPU.aluIn1\[25\] VGND VGND VPWR VPWR _04468_ sky130_fd_sc_hd__inv_2
X_14660__768 clknet_1_1__leaf__02681_ VGND VGND VPWR VPWR net800 sky130_fd_sc_hd__inv_2
Xhold1087 CPU.registerFile\[6\]\[25\] VGND VGND VPWR VPWR net2328 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1098 CPU.registerFile\[2\]\[9\] VGND VGND VPWR VPWR net2339 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_205 _07914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_216 _08397_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_227 clknet_1_0__leaf__02708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_238 _02887_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08679_ CPU.aluIn1\[11\] VGND VGND VPWR VPWR _04399_ sky130_fd_sc_hd__inv_2
XANTENNA_249 _03497_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10710_ _06048_ VGND VGND VPWR VPWR _02145_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11690_ mapped_spi_ram.rcv_data\[15\] _06588_ VGND VGND VPWR VPWR _06598_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10641_ mapped_spi_flash.rcv_data\[3\] _05994_ VGND VGND VPWR VPWR _06005_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13360_ CPU.registerFile\[21\]\[13\] _07281_ _07521_ CPU.registerFile\[17\]\[13\]
+ _07285_ VGND VGND VPWR VPWR _07790_ sky130_fd_sc_hd__o221a_1
X_10572_ mapped_spi_flash.rcv_bitcount\[3\] _05963_ VGND VGND VPWR VPWR _05964_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12311_ net2522 _06968_ _06861_ VGND VGND VPWR VPWR _06969_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13291_ _07398_ _07722_ VGND VGND VPWR VPWR _07723_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12242_ CPU.aluReg\[19\] CPU.aluReg\[17\] _06906_ VGND VGND VPWR VPWR _06916_ sky130_fd_sc_hd__mux2_1
X_12173_ CPU.aluShamt\[4\] _04286_ _06854_ VGND VGND VPWR VPWR _06864_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_31_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11124_ _06268_ VGND VGND VPWR VPWR _01951_ sky130_fd_sc_hd__clkbuf_1
X_16981_ clknet_leaf_21_clk _01307_ VGND VGND VPWR VPWR CPU.rs2\[12\] sky130_fd_sc_hd__dfxtp_1
X_11055_ _06231_ VGND VGND VPWR VPWR _01983_ sky130_fd_sc_hd__clkbuf_1
X_15932_ _03414_ _03415_ _08400_ VGND VGND VPWR VPWR _03416_ sky130_fd_sc_hd__mux2_1
X_10006_ _05597_ VGND VGND VPWR VPWR _02413_ sky130_fd_sc_hd__clkbuf_1
X_15863_ _02885_ _03346_ _03347_ _03348_ _03054_ VGND VGND VPWR VPWR _03349_ sky130_fd_sc_hd__a221o_1
X_15166__1192 clknet_1_1__leaf__02747_ VGND VGND VPWR VPWR net1224 sky130_fd_sc_hd__inv_2
X_17602_ net791 _01890_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_15794_ _02797_ _03278_ _03279_ _03281_ _03054_ VGND VGND VPWR VPWR _03282_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_35_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17533_ net722 _01821_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_106_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11957_ _06745_ VGND VGND VPWR VPWR _01592_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_106_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10908_ _06153_ VGND VGND VPWR VPWR _02052_ sky130_fd_sc_hd__clkbuf_1
X_17464_ net653 _01752_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11888_ net2523 _05735_ _06674_ VGND VGND VPWR VPWR _06709_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16415_ _02924_ _03882_ _03883_ _03884_ _02782_ VGND VGND VPWR VPWR _03885_ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13627_ _07397_ _08033_ _08048_ _08015_ VGND VGND VPWR VPWR _08049_ sky130_fd_sc_hd__a211o_1
XFILLER_0_157_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10839_ _06116_ VGND VGND VPWR VPWR _02084_ sky130_fd_sc_hd__clkbuf_1
X_17395_ net584 _01683_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_17_Left_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16346_ _03812_ _03814_ _03817_ _02965_ VGND VGND VPWR VPWR _03818_ sky130_fd_sc_hd__o22a_1
X_13558_ CPU.registerFile\[27\]\[19\] _07363_ _07981_ VGND VGND VPWR VPWR _07982_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_42_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_132_Right_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12509_ net2103 _05721_ _07071_ VGND VGND VPWR VPWR _07076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16277_ CPU.registerFile\[20\]\[25\] CPU.registerFile\[22\]\[25\] _05439_ VGND VGND
+ VPWR VPWR _03751_ sky130_fd_sc_hd__mux2_1
X_13489_ CPU.registerFile\[2\]\[17\] CPU.registerFile\[3\]\[17\] _07311_ VGND VGND
+ VPWR VPWR _07915_ sky130_fd_sc_hd__mux2_1
X_16926__6 clknet_1_1__leaf__07220_ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__inv_2
X_18016_ net1189 _02296_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_26_Left_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09720_ _05275_ _05213_ _05409_ VGND VGND VPWR VPWR _05410_ sky130_fd_sc_hd__o21a_1
XFILLER_0_129_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_143_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09651_ _04879_ _04867_ VGND VGND VPWR VPWR _05344_ sky130_fd_sc_hd__or2b_1
X_08602_ CPU.aluIn1\[11\] _04320_ VGND VGND VPWR VPWR _04322_ sky130_fd_sc_hd__nor2_1
X_09582_ _05275_ _05112_ VGND VGND VPWR VPWR _05277_ sky130_fd_sc_hd__nand2_2
X_08533_ _04251_ CPU.aluIn1\[17\] VGND VGND VPWR VPWR _04253_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_46_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_35_Left_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_154_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09016_ _04732_ VGND VGND VPWR VPWR _02578_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold140 mapped_spi_ram.cmd_addr\[8\] VGND VGND VPWR VPWR net1381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 mapped_spi_ram.cmd_addr\[6\] VGND VGND VPWR VPWR net1392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 CPU.cycles\[11\] VGND VGND VPWR VPWR net1403 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold173 mapped_spi_flash.rcv_data\[21\] VGND VGND VPWR VPWR net1414 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold184 _01712_ VGND VGND VPWR VPWR net1425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 _01713_ VGND VGND VPWR VPWR net1436 sky130_fd_sc_hd__dlygate4sd3_1
X_09918_ _05358_ VGND VGND VPWR VPWR _05547_ sky130_fd_sc_hd__clkbuf_8
X_09849_ _05500_ VGND VGND VPWR VPWR _02505_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_70_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ _07288_ _07295_ _07299_ _07301_ _07302_ VGND VGND VPWR VPWR _07303_ sky130_fd_sc_hd__a221o_1
XFILLER_0_69_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16635__80 clknet_1_1__leaf__03988_ VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__inv_2
X_11811_ _06668_ VGND VGND VPWR VPWR _01661_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_1_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _07233_ _05336_ VGND VGND VPWR VPWR _07234_ sky130_fd_sc_hd__nand2_2
XFILLER_0_95_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11742_ net1518 _06627_ _06629_ net13 VGND VGND VPWR VPWR _01692_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16650__94 clknet_1_1__leaf__03989_ VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__inv_2
XFILLER_0_139_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11673_ _06576_ VGND VGND VPWR VPWR _06588_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_48_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16200_ CPU.registerFile\[20\]\[23\] _02854_ _02819_ VGND VGND VPWR VPWR _03676_
+ sky130_fd_sc_hd__a21o_1
X_13412_ CPU.registerFile\[21\]\[15\] _07772_ _07773_ CPU.registerFile\[17\]\[15\]
+ _07839_ VGND VGND VPWR VPWR _07840_ sky130_fd_sc_hd__o221a_1
X_17180_ clknet_leaf_12_clk _01468_ VGND VGND VPWR VPWR CPU.Bimm\[3\] sky130_fd_sc_hd__dfxtp_1
X_10624_ _05967_ VGND VGND VPWR VPWR _05996_ sky130_fd_sc_hd__buf_2
XFILLER_0_24_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_742 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16131_ CPU.registerFile\[28\]\[21\] _03064_ VGND VGND VPWR VPWR _03609_ sky130_fd_sc_hd__or2_1
X_13343_ _07237_ VGND VGND VPWR VPWR _07773_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_40_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10555_ _05820_ _05950_ VGND VGND VPWR VPWR _05952_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_77_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16062_ CPU.registerFile\[19\]\[19\] CPU.registerFile\[17\]\[19\] _03025_ VGND VGND
+ VPWR VPWR _03542_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13274_ CPU.registerFile\[18\]\[11\] CPU.registerFile\[22\]\[11\] _07457_ VGND VGND
+ VPWR VPWR _07706_ sky130_fd_sc_hd__mux2_1
X_10486_ _05852_ _05895_ VGND VGND VPWR VPWR _05896_ sky130_fd_sc_hd__nor2_1
X_12225_ CPU.aluReg\[23\] CPU.aluReg\[21\] _06871_ VGND VGND VPWR VPWR _06903_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12156_ _05402_ net1736 _06841_ VGND VGND VPWR VPWR _06851_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11107_ _06259_ VGND VGND VPWR VPWR _01959_ sky130_fd_sc_hd__clkbuf_1
X_16964_ net259 _01290_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_12087_ _06814_ VGND VGND VPWR VPWR _01530_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_108_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15915_ CPU.registerFile\[14\]\[15\] CPU.registerFile\[10\]\[15\] _02849_ VGND VGND
+ VPWR VPWR _03399_ sky130_fd_sc_hd__mux2_1
X_11038_ _06222_ VGND VGND VPWR VPWR _01991_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_108_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16895_ _06030_ net1520 VGND VGND VPWR VPWR _02634_ sky130_fd_sc_hd__nor2_1
X_14643__752 clknet_1_0__leaf__02680_ VGND VGND VPWR VPWR net784 sky130_fd_sc_hd__inv_2
X_15846_ CPU.aluIn1\[12\] _03081_ _03332_ _03080_ VGND VGND VPWR VPWR _02426_ sky130_fd_sc_hd__o211a_1
X_15777_ CPU.registerFile\[14\]\[11\] CPU.registerFile\[10\]\[11\] _03082_ VGND VGND
+ VPWR VPWR _03265_ sky130_fd_sc_hd__mux2_1
X_12989_ _07238_ VGND VGND VPWR VPWR _07429_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_121_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17516_ net705 _01804_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17447_ net636 _01735_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14041__318 clknet_1_1__leaf__08364_ VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__inv_2
X_17378_ net567 _01666_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16329_ CPU.registerFile\[11\]\[27\] _02777_ VGND VGND VPWR VPWR _03801_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14726__827 clknet_1_1__leaf__02688_ VGND VGND VPWR VPWR net859 sky130_fd_sc_hd__inv_2
XFILLER_0_4_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09703_ _04410_ _04414_ VGND VGND VPWR VPWR _05394_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09634_ _04881_ _04865_ VGND VGND VPWR VPWR _05328_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09565_ _04425_ _05260_ VGND VGND VPWR VPWR _05261_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_43_Left_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08516_ CPU.aluIn1\[24\] _04235_ VGND VGND VPWR VPWR _04236_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09496_ _04889_ _05194_ VGND VGND VPWR VPWR _05195_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_156_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14772__869 clknet_1_1__leaf__02692_ VGND VGND VPWR VPWR net901 sky130_fd_sc_hd__inv_2
XFILLER_0_73_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_550 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16532__199 clknet_1_0__leaf__03964_ VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__inv_2
X_15165__1191 clknet_1_1__leaf__02747_ VGND VGND VPWR VPWR net1223 sky130_fd_sc_hd__inv_2
XFILLER_0_144_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10340_ _05791_ VGND VGND VPWR VPWR _02258_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_52_Left_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10271_ _05754_ VGND VGND VPWR VPWR _02305_ sky130_fd_sc_hd__clkbuf_1
X_12010_ _05273_ net2380 _06769_ VGND VGND VPWR VPWR _06774_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14365__502 clknet_1_0__leaf__02652_ VGND VGND VPWR VPWR net534 sky130_fd_sc_hd__inv_2
X_15700_ _02757_ _03167_ _03176_ _03190_ _02846_ VGND VGND VPWR VPWR _03191_ sky130_fd_sc_hd__a311o_2
X_12912_ _07351_ _07353_ VGND VGND VPWR VPWR _07354_ sky130_fd_sc_hd__or2_1
X_16680_ _08457_ _04005_ _04007_ _04008_ VGND VGND VPWR VPWR _04009_ sky130_fd_sc_hd__a31o_1
X_13892_ _08303_ _08304_ _07315_ VGND VGND VPWR VPWR _08305_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_61_Left_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15631_ _02760_ VGND VGND VPWR VPWR _03123_ sky130_fd_sc_hd__clkbuf_2
X_12843_ CPU.registerFile\[9\]\[0\] _07283_ _07284_ _07272_ _07285_ VGND VGND VPWR
+ VPWR _07286_ sky130_fd_sc_hd__o221a_1
XFILLER_0_158_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_87_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18350_ clknet_leaf_1_clk _02630_ VGND VGND VPWR VPWR per_uart.uart0.rx_bitcount\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_15562_ _03049_ _03055_ _02810_ VGND VGND VPWR VPWR _03056_ sky130_fd_sc_hd__a21o_1
X_17301_ net490 _01589_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11725_ net1308 mapped_spi_ram.div_counter\[1\] VGND VGND VPWR VPWR _06617_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_25_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18281_ net114 _02561_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_15493_ CPU.registerFile\[22\]\[3\] CPU.registerFile\[23\]\[3\] _02829_ VGND VGND
+ VPWR VPWR _02989_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17232_ net422 _01520_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[25\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03970_ _03970_ VGND VGND VPWR VPWR clknet_0__03970_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_154_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11656_ mapped_spi_ram.rcv_data\[30\] _06577_ VGND VGND VPWR VPWR _06579_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17163_ net387 _01451_ VGND VGND VPWR VPWR CPU.aluReg\[27\] sky130_fd_sc_hd__dfxtp_1
X_10607_ net1458 _05983_ _05986_ _05980_ VGND VGND VPWR VPWR _02185_ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11587_ net1375 _06517_ _06509_ _06529_ VGND VGND VPWR VPWR _06530_ sky130_fd_sc_hd__a211o_1
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16114_ CPU.registerFile\[28\]\[20\] CPU.registerFile\[24\]\[20\] _02761_ VGND VGND
+ VPWR VPWR _03593_ sky130_fd_sc_hd__mux2_1
X_13326_ CPU.registerFile\[13\]\[12\] _07281_ _07521_ CPU.registerFile\[9\]\[12\]
+ _07285_ VGND VGND VPWR VPWR _07757_ sky130_fd_sc_hd__o221a_1
XFILLER_0_40_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17094_ net352 _01416_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__02752_ clknet_0__02752_ VGND VGND VPWR VPWR clknet_1_1__leaf__02752_
+ sky130_fd_sc_hd__clkbuf_16
X_10538_ net1442 _05892_ _05938_ _05936_ VGND VGND VPWR VPWR _02206_ sky130_fd_sc_hd__o211a_1
Xhold909 CPU.registerFile\[21\]\[12\] VGND VGND VPWR VPWR net2150 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16045_ CPU.registerFile\[18\]\[18\] _03068_ _03069_ CPU.registerFile\[19\]\[18\]
+ _03074_ VGND VGND VPWR VPWR _03526_ sky130_fd_sc_hd__o221a_1
X_13257_ CPU.registerFile\[29\]\[10\] _07414_ _07326_ CPU.registerFile\[25\]\[10\]
+ _07489_ VGND VGND VPWR VPWR _07690_ sky130_fd_sc_hd__o221a_1
X_10469_ _04507_ _04551_ _04552_ _04629_ VGND VGND VPWR VPWR _05881_ sky130_fd_sc_hd__a31o_1
XFILLER_0_122_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__02683_ clknet_0__02683_ VGND VGND VPWR VPWR clknet_1_1__leaf__02683_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_122_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12208_ CPU.aluIn1\[26\] _06889_ _06865_ VGND VGND VPWR VPWR _06890_ sky130_fd_sc_hd__mux2_1
X_13188_ CPU.registerFile\[11\]\[8\] _07619_ _07622_ VGND VGND VPWR VPWR _07623_ sky130_fd_sc_hd__o21a_1
X_12139_ _06842_ VGND VGND VPWR VPWR _01506_ sky130_fd_sc_hd__clkbuf_1
X_17996_ clknet_leaf_8_clk _02280_ VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[10\]
+ sky130_fd_sc_hd__dfxtp_1
X_16947_ net242 _01273_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_16878_ per_uart.uart0.rx_count16\[3\] per_uart.uart0.rx_count16\[2\] _04156_ VGND
+ VGND VPWR VPWR _04162_ sky130_fd_sc_hd__nand3_1
X_15829_ _03311_ _03315_ _03138_ VGND VGND VPWR VPWR _03316_ sky130_fd_sc_hd__a21o_1
X_09350_ _04800_ _05055_ VGND VGND VPWR VPWR _05056_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09281_ CPU.Iimm\[0\] _04812_ _04989_ CPU.cycles\[20\] VGND VGND VPWR VPWR _04990_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_151_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload60 clknet_1_1__leaf__02695_ VGND VGND VPWR VPWR clkload60/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload71 clknet_1_1__leaf__02664_ VGND VGND VPWR VPWR clkload71/X sky130_fd_sc_hd__clkbuf_8
Xclkload82 clknet_1_1__leaf__02662_ VGND VGND VPWR VPWR clkload82/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_141_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload93 clknet_1_0__leaf__08466_ VGND VGND VPWR VPWR clkload93/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_100_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14314__456 clknet_1_1__leaf__08464_ VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__inv_2
X_08996_ _04713_ VGND VGND VPWR VPWR _04714_ sky130_fd_sc_hd__buf_8
X_13952__238 clknet_1_0__leaf__07226_ VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_149_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09617_ _04218_ _04621_ VGND VGND VPWR VPWR _05311_ sky130_fd_sc_hd__nand2_1
X_09548_ _04426_ _05244_ VGND VGND VPWR VPWR _05245_ sky130_fd_sc_hd__xor2_1
XFILLER_0_93_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09479_ _04974_ _05175_ _05178_ VGND VGND VPWR VPWR _05179_ sky130_fd_sc_hd__o21ai_2
X_14360__498 clknet_1_0__leaf__08468_ VGND VGND VPWR VPWR net530 sky130_fd_sc_hd__inv_2
XFILLER_0_148_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11510_ CPU.mem_rstrb _05068_ _06468_ net1336 VGND VGND VPWR VPWR _06476_ sky130_fd_sc_hd__and4b_1
XFILLER_0_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12490_ net1753 _05702_ _07060_ VGND VGND VPWR VPWR _07066_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11441_ _05497_ CPU.registerFile\[25\]\[28\] _06433_ VGND VGND VPWR VPWR _06437_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14160_ CPU.Iimm\[3\] _07397_ _08413_ VGND VGND VPWR VPWR _08417_ sky130_fd_sc_hd__mux2_1
X_11372_ _06400_ VGND VGND VPWR VPWR _01835_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13111_ CPU.registerFile\[8\]\[6\] CPU.registerFile\[12\]\[6\] _07314_ VGND VGND
+ VPWR VPWR _07548_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10323_ _05782_ VGND VGND VPWR VPWR _02266_ sky130_fd_sc_hd__clkbuf_1
X_14091_ _04650_ _07128_ VGND VGND VPWR VPWR _08372_ sky130_fd_sc_hd__nor2_1
X_13042_ CPU.registerFile\[30\]\[4\] CPU.registerFile\[26\]\[4\] _07480_ VGND VGND
+ VPWR VPWR _07481_ sky130_fd_sc_hd__mux2_1
X_10254_ _05745_ VGND VGND VPWR VPWR _02313_ sky130_fd_sc_hd__clkbuf_1
X_14709__811 clknet_1_0__leaf__02687_ VGND VGND VPWR VPWR net843 sky130_fd_sc_hd__inv_2
X_17850_ net1039 _02134_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_10185_ _05699_ VGND VGND VPWR VPWR _02336_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14289__433 clknet_1_1__leaf__08462_ VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__inv_2
XFILLER_0_100_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14070__344 clknet_1_1__leaf__08367_ VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__inv_2
X_16801_ _04106_ _04110_ _05815_ VGND VGND VPWR VPWR _02603_ sky130_fd_sc_hd__a21oi_1
X_17781_ net970 _02065_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_16732_ _04052_ _05155_ _04006_ VGND VGND VPWR VPWR _04053_ sky130_fd_sc_hd__or3b_1
X_13944_ per_uart.uart0.enable16_counter\[15\] _07193_ VGND VGND VPWR VPWR _08355_
+ sky130_fd_sc_hd__nor2_2
X_16663_ _05288_ _08454_ _05390_ VGND VGND VPWR VPWR _03994_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_85_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13875_ CPU.registerFile\[31\]\[29\] _07556_ _07557_ CPU.registerFile\[27\]\[29\]
+ _08288_ VGND VGND VPWR VPWR _08289_ sky130_fd_sc_hd__o221a_1
XFILLER_0_158_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12826_ _07254_ _07259_ _07267_ _07268_ VGND VGND VPWR VPWR _07269_ sky130_fd_sc_hd__o211a_1
X_15614_ CPU.registerFile\[22\]\[6\] CPU.registerFile\[23\]\[6\] _02829_ VGND VGND
+ VPWR VPWR _03107_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18333_ clknet_leaf_6_clk _02613_ VGND VGND VPWR VPWR per_uart.uart0.tx_bitcount\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_15545_ CPU.registerFile\[8\]\[5\] _02763_ _02764_ _03038_ VGND VGND VPWR VPWR _03039_
+ sky130_fd_sc_hd__o211a_1
X_12757_ clknet_2_0__leaf_clk VGND VGND VPWR VPWR _07222_ sky130_fd_sc_hd__buf_1
XFILLER_0_155_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14755__853 clknet_1_0__leaf__02691_ VGND VGND VPWR VPWR net885 sky130_fd_sc_hd__inv_2
X_11708_ net2378 _06603_ _06608_ _06607_ VGND VGND VPWR VPWR _01703_ sky130_fd_sc_hd__o211a_1
X_15476_ CPU.registerFile\[27\]\[3\] CPU.registerFile\[31\]\[3\] _02852_ VGND VGND
+ VPWR VPWR _02972_ sky130_fd_sc_hd__mux2_1
X_18264_ clknet_leaf_2_clk _02544_ VGND VGND VPWR VPWR per_uart.uart0.rxd_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_12688_ CPU.cycles\[28\] _07170_ net1421 VGND VGND VPWR VPWR _07173_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16515__183 clknet_1_0__leaf__03963_ VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__inv_2
X_17215_ net405 _01503_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11639_ net1494 _06562_ _06565_ _06492_ VGND VGND VPWR VPWR _01729_ sky130_fd_sc_hd__a22o_1
X_18195_ net226 _02475_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_15005__1079 clknet_1_0__leaf__02715_ VGND VGND VPWR VPWR net1111 sky130_fd_sc_hd__inv_2
XFILLER_0_142_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17146_ net370 _01434_ VGND VGND VPWR VPWR CPU.aluReg\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold706 CPU.registerFile\[3\]\[15\] VGND VGND VPWR VPWR net1947 sky130_fd_sc_hd__dlygate4sd3_1
Xhold717 CPU.registerFile\[1\]\[28\] VGND VGND VPWR VPWR net1958 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold728 CPU.registerFile\[23\]\[21\] VGND VGND VPWR VPWR net1969 sky130_fd_sc_hd__dlygate4sd3_1
X_13309_ CPU.registerFile\[23\]\[12\] _07244_ _07239_ CPU.registerFile\[19\]\[12\]
+ _07739_ VGND VGND VPWR VPWR _07740_ sky130_fd_sc_hd__o221a_1
X_17077_ net335 _01399_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[7\] sky130_fd_sc_hd__dfxtp_1
Xhold739 CPU.registerFile\[30\]\[20\] VGND VGND VPWR VPWR net1980 sky130_fd_sc_hd__dlygate4sd3_1
X_16028_ CPU.registerFile\[24\]\[18\] _03130_ _02780_ _03508_ VGND VGND VPWR VPWR
+ _03509_ sky130_fd_sc_hd__o211a_1
Xclkbuf_1_1__f__02666_ clknet_0__02666_ VGND VGND VPWR VPWR clknet_1_1__leaf__02666_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_110_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08850_ CPU.aluIn1\[19\] CPU.aluIn1\[18\] _04495_ VGND VGND VPWR VPWR _04570_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_0__02697_ _02697_ VGND VGND VPWR VPWR clknet_0__02697_ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_0__07224_ _07224_ VGND VGND VPWR VPWR clknet_0__07224_ sky130_fd_sc_hd__clkbuf_16
X_08781_ _04500_ _04291_ _04292_ _04294_ VGND VGND VPWR VPWR _04501_ sky130_fd_sc_hd__and4_1
XFILLER_0_46_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17979_ net1167 _02263_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_15164__1190 clknet_1_0__leaf__02747_ VGND VGND VPWR VPWR net1222 sky130_fd_sc_hd__inv_2
XFILLER_0_79_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09402_ _04331_ _04211_ _04219_ CPU.aluReg\[15\] _05105_ VGND VGND VPWR VPWR _05106_
+ sky130_fd_sc_hd__a221o_1
X_14838__928 clknet_1_0__leaf__02699_ VGND VGND VPWR VPWR net960 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_9_Left_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09333_ _05033_ _05039_ _04773_ VGND VGND VPWR VPWR _05040_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09264_ _04817_ VGND VGND VPWR VPWR _04974_ sky130_fd_sc_hd__buf_4
XFILLER_0_56_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09195_ _04827_ _04906_ VGND VGND VPWR VPWR _04907_ sky130_fd_sc_hd__and2_1
XFILLER_0_145_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15221__131 clknet_1_1__leaf__02753_ VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__inv_2
XFILLER_0_87_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08979_ _04697_ VGND VGND VPWR VPWR _02580_ sky130_fd_sc_hd__clkbuf_1
Xhold77 mapped_spi_ram.cmd_addr\[30\] VGND VGND VPWR VPWR net1318 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ _06763_ VGND VGND VPWR VPWR _01577_ sky130_fd_sc_hd__clkbuf_1
Xhold88 mapped_spi_flash.state\[0\] VGND VGND VPWR VPWR net1329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 _02730_ VGND VGND VPWR VPWR net1340 sky130_fd_sc_hd__dlygate4sd3_1
X_10941_ net1554 _05723_ _06165_ VGND VGND VPWR VPWR _06171_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__02755_ clknet_0__02755_ VGND VGND VPWR VPWR clknet_1_0__leaf__02755_
+ sky130_fd_sc_hd__clkbuf_16
X_13660_ CPU.registerFile\[30\]\[23\] _07987_ VGND VGND VPWR VPWR _08080_ sky130_fd_sc_hd__or2_1
X_10872_ net2422 _05723_ _06128_ VGND VGND VPWR VPWR _06134_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__02686_ clknet_0__02686_ VGND VGND VPWR VPWR clknet_1_0__leaf__02686_
+ sky130_fd_sc_hd__clkbuf_16
X_12611_ _05816_ net1498 VGND VGND VPWR VPWR _07129_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13591_ _07334_ _08003_ _08006_ _08013_ _07766_ VGND VGND VPWR VPWR _08014_ sky130_fd_sc_hd__o311a_1
XFILLER_0_66_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14477__603 clknet_1_0__leaf__02663_ VGND VGND VPWR VPWR net635 sky130_fd_sc_hd__inv_2
XFILLER_0_137_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15330_ _02828_ VGND VGND VPWR VPWR _02829_ sky130_fd_sc_hd__buf_4
X_12542_ _07093_ VGND VGND VPWR VPWR _01287_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_80_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15261_ _05048_ VGND VGND VPWR VPWR _02760_ sky130_fd_sc_hd__buf_4
XFILLER_0_151_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12473_ net2291 _05685_ _07049_ VGND VGND VPWR VPWR _07057_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_412 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17000_ clknet_leaf_21_clk _01326_ VGND VGND VPWR VPWR CPU.rs2\[31\] sky130_fd_sc_hd__dfxtp_1
X_11424_ _06427_ VGND VGND VPWR VPWR _01810_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_8 _02819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14143_ CPU.Jimm\[17\] _08405_ _08387_ VGND VGND VPWR VPWR _08406_ sky130_fd_sc_hd__mux2_1
X_11355_ _06390_ VGND VGND VPWR VPWR _01842_ sky130_fd_sc_hd__clkbuf_1
X_10306_ _05772_ VGND VGND VPWR VPWR _02288_ sky130_fd_sc_hd__clkbuf_1
X_11286_ CPU.registerFile\[9\]\[4\] _05727_ _06346_ VGND VGND VPWR VPWR _06354_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13025_ _07369_ _07461_ _07463_ _07231_ VGND VGND VPWR VPWR _07464_ sky130_fd_sc_hd__a211o_1
X_17902_ net1091 _02186_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_111_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10237_ _05734_ VGND VGND VPWR VPWR _02319_ sky130_fd_sc_hd__clkbuf_1
X_17482__28 VGND VGND VPWR VPWR _17482__28/HI net28 sky130_fd_sc_hd__conb_1
X_17833_ net1022 _02117_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_10168_ net2142 _05687_ _05671_ VGND VGND VPWR VPWR _05688_ sky130_fd_sc_hd__mux2_1
X_17764_ net953 _02048_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10099_ net1631 _05027_ _05644_ VGND VGND VPWR VPWR _05647_ sky130_fd_sc_hd__mux2_1
X_16715_ _03991_ net2427 VGND VGND VPWR VPWR _04038_ sky130_fd_sc_hd__nand2_1
X_13927_ _07360_ _08328_ _08331_ _08338_ VGND VGND VPWR VPWR _08339_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17695_ net884 _01983_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_14919__1001 clknet_1_1__leaf__02707_ VGND VGND VPWR VPWR net1033 sky130_fd_sc_hd__inv_2
X_13858_ CPU.registerFile\[1\]\[29\] _07387_ _08271_ _07379_ VGND VGND VPWR VPWR _08272_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_85_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12809_ _05308_ VGND VGND VPWR VPWR _07252_ sky130_fd_sc_hd__buf_4
X_14343__482 clknet_1_0__leaf__08467_ VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__inv_2
X_16577_ clknet_1_1__leaf__07219_ VGND VGND VPWR VPWR _03969_ sky130_fd_sc_hd__buf_1
XFILLER_0_128_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13789_ CPU.registerFile\[6\]\[27\] CPU.registerFile\[7\]\[27\] _07641_ VGND VGND
+ VPWR VPWR _08205_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18316_ clknet_leaf_16_clk _02596_ VGND VGND VPWR VPWR CPU.PC\[16\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_57_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15528_ CPU.registerFile\[21\]\[4\] CPU.registerFile\[23\]\[4\] _02769_ VGND VGND
+ VPWR VPWR _03023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13981__264 clknet_1_0__leaf__08358_ VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18247_ net88 _02527_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15459_ _02949_ _02952_ _02955_ VGND VGND VPWR VPWR _02956_ sky130_fd_sc_hd__or3_2
X_18178_ net209 _02458_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold503 CPU.registerFile\[9\]\[31\] VGND VGND VPWR VPWR net1744 sky130_fd_sc_hd__dlygate4sd3_1
X_17129_ clknet_leaf_22_clk _00032_ VGND VGND VPWR VPWR CPU.cycles\[25\] sky130_fd_sc_hd__dfxtp_1
Xhold514 mapped_spi_ram.rcv_bitcount\[5\] VGND VGND VPWR VPWR net1755 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold525 CPU.registerFile\[20\]\[14\] VGND VGND VPWR VPWR net1766 sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 CPU.registerFile\[16\]\[6\] VGND VGND VPWR VPWR net1777 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold547 CPU.registerFile\[29\]\[28\] VGND VGND VPWR VPWR net1788 sky130_fd_sc_hd__dlygate4sd3_1
X_09951_ _05567_ VGND VGND VPWR VPWR _02470_ sky130_fd_sc_hd__clkbuf_1
Xhold558 CPU.registerFile\[26\]\[3\] VGND VGND VPWR VPWR net1799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 CPU.registerFile\[21\]\[15\] VGND VGND VPWR VPWR net1810 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__02718_ clknet_0__02718_ VGND VGND VPWR VPWR clknet_1_1__leaf__02718_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_21_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08902_ net15 _04619_ _04621_ VGND VGND VPWR VPWR _04622_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__02749_ _02749_ VGND VGND VPWR VPWR clknet_0__02749_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_148_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09882_ _05522_ net2406 _05512_ VGND VGND VPWR VPWR _05523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08833_ _04552_ _04551_ VGND VGND VPWR VPWR _04553_ sky130_fd_sc_hd__or2_4
XFILLER_0_148_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1203 CPU.registerFile\[23\]\[7\] VGND VGND VPWR VPWR net2444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1214 CPU.registerFile\[20\]\[17\] VGND VGND VPWR VPWR net2455 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1225 CPU.registerFile\[10\]\[6\] VGND VGND VPWR VPWR net2466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_146_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1236 CPU.registerFile\[25\]\[14\] VGND VGND VPWR VPWR net2477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1247 CPU.registerFile\[8\]\[2\] VGND VGND VPWR VPWR net2488 sky130_fd_sc_hd__dlygate4sd3_1
X_08764_ CPU.Jimm\[13\] CPU.Jimm\[12\] VGND VGND VPWR VPWR _04484_ sky130_fd_sc_hd__or2_4
Xhold1258 CPU.registerFile\[10\]\[3\] VGND VGND VPWR VPWR net2499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 CPU.registerFile\[8\]\[9\] VGND VGND VPWR VPWR net2510 sky130_fd_sc_hd__dlygate4sd3_1
X_08695_ _04288_ CPU.aluIn1\[2\] VGND VGND VPWR VPWR _04415_ sky130_fd_sc_hd__xor2_4
XANTENNA_409 _04659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14426__557 clknet_1_1__leaf__02658_ VGND VGND VPWR VPWR net589 sky130_fd_sc_hd__inv_2
XFILLER_0_79_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_146_Right_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09316_ _04927_ _05023_ VGND VGND VPWR VPWR _05024_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09247_ _04957_ VGND VGND VPWR VPWR _04958_ sky130_fd_sc_hd__buf_4
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09178_ CPU.Bimm\[10\] _04820_ CPU.PC\[10\] VGND VGND VPWR VPWR _04890_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_478 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput12 net12 VGND VGND VPWR VPWR spi_mosi_ram sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14472__599 clknet_1_1__leaf__02662_ VGND VGND VPWR VPWR net631 sky130_fd_sc_hd__inv_2
X_11140_ net2510 _05717_ _06274_ VGND VGND VPWR VPWR _06277_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11071_ net1912 _05717_ _06237_ VGND VGND VPWR VPWR _06240_ sky130_fd_sc_hd__mux2_1
X_10022_ _05605_ VGND VGND VPWR VPWR _02405_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15004__1078 clknet_1_0__leaf__02715_ VGND VGND VPWR VPWR net1110 sky130_fd_sc_hd__inv_2
X_11973_ _06754_ VGND VGND VPWR VPWR _01585_ sky130_fd_sc_hd__clkbuf_1
X_16500_ clknet_1_0__leaf__02749_ VGND VGND VPWR VPWR _03962_ sky130_fd_sc_hd__buf_1
X_10924_ net1775 _05706_ _06154_ VGND VGND VPWR VPWR _06162_ sky130_fd_sc_hd__mux2_1
X_13712_ CPU.registerFile\[13\]\[24\] _07361_ _08130_ _07417_ _07554_ VGND VGND VPWR
+ VPWR _08131_ sky130_fd_sc_hd__o221a_1
XFILLER_0_85_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17480_ net669 net26 VGND VGND VPWR VPWR mapped_spi_flash.div_counter\[3\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_113_Right_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16431_ CPU.registerFile\[14\]\[30\] CPU.registerFile\[10\]\[30\] _02761_ VGND VGND
+ VPWR VPWR _03900_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10855_ CPU.registerFile\[2\]\[14\] _05706_ _06117_ VGND VGND VPWR VPWR _06125_ sky130_fd_sc_hd__mux2_1
X_13643_ _07646_ _08053_ _08056_ _08063_ VGND VGND VPWR VPWR _08064_ sky130_fd_sc_hd__a31o_1
XFILLER_0_67_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__02669_ clknet_0__02669_ VGND VGND VPWR VPWR clknet_1_0__leaf__02669_
+ sky130_fd_sc_hd__clkbuf_16
X_16362_ _02786_ _03830_ _03832_ _03019_ VGND VGND VPWR VPWR _03833_ sky130_fd_sc_hd__a211o_1
X_13574_ CPU.registerFile\[21\]\[20\] _07244_ _07429_ CPU.registerFile\[17\]\[20\]
+ _07349_ VGND VGND VPWR VPWR _07997_ sky130_fd_sc_hd__o221a_1
XFILLER_0_39_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10786_ _06088_ VGND VGND VPWR VPWR _02109_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18101_ net164 _02381_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_12525_ _04662_ _06141_ VGND VGND VPWR VPWR _07084_ sky130_fd_sc_hd__nor2_2
X_15313_ _02758_ VGND VGND VPWR VPWR _02812_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_30_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16293_ _03764_ _03765_ _02856_ VGND VGND VPWR VPWR _03766_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18032_ net1205 _02312_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_12456_ _07047_ VGND VGND VPWR VPWR _01360_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11407_ _06418_ VGND VGND VPWR VPWR _01818_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12387_ _05448_ net1919 _06976_ VGND VGND VPWR VPWR _07011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14867__954 clknet_1_0__leaf__02702_ VGND VGND VPWR VPWR net986 sky130_fd_sc_hd__inv_2
X_14126_ _08392_ VGND VGND VPWR VPWR _01471_ sky130_fd_sc_hd__clkbuf_1
X_11338_ _06381_ VGND VGND VPWR VPWR _01850_ sky130_fd_sc_hd__clkbuf_1
X_11269_ CPU.registerFile\[9\]\[12\] _05710_ _06335_ VGND VGND VPWR VPWR _06345_ sky130_fd_sc_hd__mux2_1
X_13008_ CPU.registerFile\[30\]\[3\] CPU.registerFile\[26\]\[3\] _07292_ VGND VGND
+ VPWR VPWR _07448_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17816_ net1005 _02100_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_128_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17747_ net936 _02031_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08480_ _04199_ VGND VGND VPWR VPWR _04200_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_141_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17678_ net867 _01966_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_141_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09101_ CPU.Iimm\[3\] _04812_ _04503_ CPU.cycles\[23\] VGND VGND VPWR VPWR _04813_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_44_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_99_Left_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_866 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09032_ _04747_ VGND VGND VPWR VPWR _04748_ sky130_fd_sc_hd__buf_2
XFILLER_0_142_220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold300 _04141_ VGND VGND VPWR VPWR net1541 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold311 per_uart.uart0.rxd_reg\[3\] VGND VGND VPWR VPWR net1552 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold322 CPU.registerFile\[6\]\[4\] VGND VGND VPWR VPWR net1563 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold333 CPU.registerFile\[5\]\[18\] VGND VGND VPWR VPWR net1574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold344 CPU.registerFile\[5\]\[8\] VGND VGND VPWR VPWR net1585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 CPU.registerFile\[30\]\[23\] VGND VGND VPWR VPWR net1596 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold366 CPU.registerFile\[6\]\[27\] VGND VGND VPWR VPWR net1607 sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 CPU.registerFile\[17\]\[23\] VGND VGND VPWR VPWR net1618 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold388 CPU.registerFile\[14\]\[23\] VGND VGND VPWR VPWR net1629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold399 CPU.registerFile\[7\]\[4\] VGND VGND VPWR VPWR net1640 sky130_fd_sc_hd__dlygate4sd3_1
X_09934_ _05489_ _05557_ VGND VGND VPWR VPWR _05558_ sky130_fd_sc_hd__nand2_2
X_09865_ _04981_ VGND VGND VPWR VPWR _05511_ sky130_fd_sc_hd__clkbuf_4
Xhold1000 CPU.registerFile\[15\]\[15\] VGND VGND VPWR VPWR net2241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1011 CPU.registerFile\[27\]\[13\] VGND VGND VPWR VPWR net2252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1022 CPU.registerFile\[12\]\[4\] VGND VGND VPWR VPWR net2263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1033 CPU.registerFile\[22\]\[6\] VGND VGND VPWR VPWR net2274 sky130_fd_sc_hd__dlygate4sd3_1
X_08816_ CPU.aluIn1\[5\] CPU.Bimm\[5\] VGND VGND VPWR VPWR _04536_ sky130_fd_sc_hd__or2_1
Xhold1044 CPU.registerFile\[26\]\[27\] VGND VGND VPWR VPWR net2285 sky130_fd_sc_hd__dlygate4sd3_1
X_09796_ net2333 _05090_ _05463_ VGND VGND VPWR VPWR _05469_ sky130_fd_sc_hd__mux2_1
Xhold1055 per_uart.uart0.tx_bitcount\[3\] VGND VGND VPWR VPWR net2296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 CPU.registerFile\[4\]\[16\] VGND VGND VPWR VPWR net2307 sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ _04465_ _04463_ _04359_ _04466_ _04353_ VGND VGND VPWR VPWR _04467_ sky130_fd_sc_hd__a2111o_1
Xhold1077 CPU.registerFile\[23\]\[22\] VGND VGND VPWR VPWR net2318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1088 CPU.registerFile\[14\]\[25\] VGND VGND VPWR VPWR net2329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1099 per_uart.uart0.tx_bitcount\[2\] VGND VGND VPWR VPWR net2340 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_206 _07914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_217 _08403_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_228 clknet_1_1__leaf__02697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_239 _02887_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08678_ _04397_ _04261_ VGND VGND VPWR VPWR _04398_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_64_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10640_ net2035 _05996_ _06004_ _05993_ VGND VGND VPWR VPWR _02170_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10571_ mapped_spi_flash.rcv_bitcount\[2\] mapped_spi_flash.rcv_bitcount\[1\] mapped_spi_flash.rcv_bitcount\[0\]
+ VGND VGND VPWR VPWR _05963_ sky130_fd_sc_hd__or3_1
XFILLER_0_64_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12310_ CPU.aluIn1\[2\] _06967_ _06859_ VGND VGND VPWR VPWR _06968_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13290_ CPU.registerFile\[30\]\[11\] CPU.registerFile\[26\]\[11\] _07399_ VGND VGND
+ VPWR VPWR _07722_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12241_ _06915_ VGND VGND VPWR VPWR _01443_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14589__704 clknet_1_0__leaf__02674_ VGND VGND VPWR VPWR net736 sky130_fd_sc_hd__inv_2
XFILLER_0_133_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12172_ CPU.aluShamt\[2\] CPU.aluShamt\[1\] CPU.aluShamt\[0\] net1542 VGND VGND VPWR
+ VPWR _06863_ sky130_fd_sc_hd__o31a_1
X_14918__1000 clknet_1_1__leaf__02707_ VGND VGND VPWR VPWR net1032 sky130_fd_sc_hd__inv_2
XFILLER_0_102_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11123_ CPU.registerFile\[8\]\[17\] _05700_ _06263_ VGND VGND VPWR VPWR _06268_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16980_ clknet_leaf_28_clk _01306_ VGND VGND VPWR VPWR CPU.rs2\[11\] sky130_fd_sc_hd__dfxtp_1
X_11054_ net2409 _05700_ _06226_ VGND VGND VPWR VPWR _06231_ sky130_fd_sc_hd__mux2_1
X_15931_ CPU.registerFile\[30\]\[15\] CPU.registerFile\[26\]\[15\] _02773_ VGND VGND
+ VPWR VPWR _03415_ sky130_fd_sc_hd__mux2_1
X_10005_ net1800 _04659_ _05596_ VGND VGND VPWR VPWR _05597_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15862_ CPU.registerFile\[25\]\[13\] _03280_ _02803_ VGND VGND VPWR VPWR _03348_
+ sky130_fd_sc_hd__o21a_1
X_17601_ net790 _01889_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_14409__541 clknet_1_0__leaf__02657_ VGND VGND VPWR VPWR net573 sky130_fd_sc_hd__inv_2
X_15793_ CPU.registerFile\[25\]\[11\] _03280_ _02803_ VGND VGND VPWR VPWR _03281_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17532_ net721 _01820_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_11956_ CPU.registerFile\[11\]\[0\] _05735_ _06710_ VGND VGND VPWR VPWR _06745_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_123_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10907_ net1710 _05689_ _06143_ VGND VGND VPWR VPWR _06153_ sky130_fd_sc_hd__mux2_1
X_17463_ net652 _01751_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[18\] sky130_fd_sc_hd__dfxtp_1
X_11887_ _06708_ VGND VGND VPWR VPWR _01625_ sky130_fd_sc_hd__clkbuf_1
X_16414_ CPU.registerFile\[13\]\[29\] _02775_ VGND VGND VPWR VPWR _03884_ sky130_fd_sc_hd__or2_1
X_10838_ net2104 _05689_ _06106_ VGND VGND VPWR VPWR _06116_ sky130_fd_sc_hd__mux2_1
X_13626_ _08040_ _08047_ _07394_ VGND VGND VPWR VPWR _08048_ sky130_fd_sc_hd__o21a_1
X_17394_ net583 _01682_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16345_ _03815_ _03816_ _02855_ VGND VGND VPWR VPWR _03817_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13557_ CPU.registerFile\[31\]\[19\] _07325_ _07980_ _07621_ _07327_ VGND VGND VPWR
+ VPWR _07981_ sky130_fd_sc_hd__o221a_1
X_10769_ _06079_ VGND VGND VPWR VPWR _02117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12508_ _07075_ VGND VGND VPWR VPWR _01336_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_229 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16276_ CPU.registerFile\[21\]\[25\] CPU.registerFile\[23\]\[25\] _05439_ VGND VGND
+ VPWR VPWR _03750_ sky130_fd_sc_hd__mux2_1
X_13488_ _07909_ _07910_ _07911_ _07913_ VGND VGND VPWR VPWR _07914_ sky130_fd_sc_hd__a22o_2
XFILLER_0_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18015_ net1188 _02295_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12439_ _05253_ net1871 _07035_ VGND VGND VPWR VPWR _07039_ sky130_fd_sc_hd__mux2_1
X_14455__583 clknet_1_0__leaf__02661_ VGND VGND VPWR VPWR net615 sky130_fd_sc_hd__inv_2
XFILLER_0_23_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14193__371 clknet_1_1__leaf__08429_ VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__inv_2
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14109_ _04291_ _05279_ _00000_ VGND VGND VPWR VPWR _08383_ sky130_fd_sc_hd__mux2_1
X_15089_ _07183_ _02731_ _02727_ VGND VGND VPWR VPWR _02274_ sky130_fd_sc_hd__a21oi_1
X_09650_ _04869_ _04878_ VGND VGND VPWR VPWR _05343_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_143_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08601_ CPU.aluIn1\[11\] _04320_ VGND VGND VPWR VPWR _04321_ sky130_fd_sc_hd__and2_1
X_09581_ _04692_ _05111_ _04636_ VGND VGND VPWR VPWR _05276_ sky130_fd_sc_hd__mux2_1
X_08532_ CPU.aluIn1\[17\] _04251_ VGND VGND VPWR VPWR _04252_ sky130_fd_sc_hd__or2b_1
XFILLER_0_77_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14620__731 clknet_1_1__leaf__02678_ VGND VGND VPWR VPWR net763 sky130_fd_sc_hd__inv_2
XFILLER_0_148_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14538__658 clknet_1_0__leaf__02669_ VGND VGND VPWR VPWR net690 sky130_fd_sc_hd__inv_2
XFILLER_0_116_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09015_ net1686 _04731_ _04668_ VGND VGND VPWR VPWR _04732_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15003__1077 clknet_1_0__leaf__02715_ VGND VGND VPWR VPWR net1109 sky130_fd_sc_hd__inv_2
XFILLER_0_14_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold130 mapped_spi_ram.cmd_addr\[15\] VGND VGND VPWR VPWR net1371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 mapped_spi_flash.cmd_addr\[7\] VGND VGND VPWR VPWR net1382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 mapped_spi_ram.cmd_addr\[24\] VGND VGND VPWR VPWR net1393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 mapped_spi_flash.rcv_data\[25\] VGND VGND VPWR VPWR net1404 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold174 _02188_ VGND VGND VPWR VPWR net1415 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold185 CPU.cycles\[31\] VGND VGND VPWR VPWR net1426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 CPU.cycles\[23\] VGND VGND VPWR VPWR net1437 sky130_fd_sc_hd__dlygate4sd3_1
X_09917_ _05546_ VGND VGND VPWR VPWR _02483_ sky130_fd_sc_hd__clkbuf_1
X_09848_ _05499_ net2438 _05491_ VGND VGND VPWR VPWR _05500_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ net2331 _04798_ _05452_ VGND VGND VPWR VPWR _05460_ sky130_fd_sc_hd__mux2_1
X_11810_ _05333_ net2348 _06661_ VGND VGND VPWR VPWR _06668_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _05282_ VGND VGND VPWR VPWR _07233_ sky130_fd_sc_hd__clkbuf_8
X_14896__980 clknet_1_0__leaf__02705_ VGND VGND VPWR VPWR net1012 sky130_fd_sc_hd__inv_2
X_11741_ _06471_ _06569_ _00008_ VGND VGND VPWR VPWR _06630_ sky130_fd_sc_hd__nor3_1
XFILLER_0_68_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11672_ net1482 _06575_ _06587_ _06581_ VGND VGND VPWR VPWR _01718_ sky130_fd_sc_hd__o211a_1
X_10623_ mapped_spi_flash.rcv_data\[11\] _05983_ _05995_ _05993_ VGND VGND VPWR VPWR
+ _02178_ sky130_fd_sc_hd__o211a_1
X_13411_ _07370_ _07838_ VGND VGND VPWR VPWR _07839_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_21_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_153_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16130_ CPU.registerFile\[30\]\[21\] CPU.registerFile\[26\]\[21\] _03247_ VGND VGND
+ VPWR VPWR _03608_ sky130_fd_sc_hd__mux2_1
X_13342_ _07234_ VGND VGND VPWR VPWR _07772_ sky130_fd_sc_hd__buf_4
XFILLER_0_107_754 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10554_ _05951_ VGND VGND VPWR VPWR _02203_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_77_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13273_ _07228_ VGND VGND VPWR VPWR _07705_ sky130_fd_sc_hd__buf_2
X_16061_ CPU.registerFile\[16\]\[19\] CPU.registerFile\[18\]\[19\] _03032_ VGND VGND
+ VPWR VPWR _03541_ sky130_fd_sc_hd__mux2_1
X_10485_ CPU.PC\[11\] _05867_ _05894_ _04629_ VGND VGND VPWR VPWR _05895_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12224_ _06902_ VGND VGND VPWR VPWR _01447_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12155_ _06850_ VGND VGND VPWR VPWR _01498_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_9_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11106_ net2443 _05683_ _06252_ VGND VGND VPWR VPWR _06259_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16963_ net258 _01289_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_12086_ _05381_ net1799 _06805_ VGND VGND VPWR VPWR _06814_ sky130_fd_sc_hd__mux2_1
X_15914_ CPU.aluIn1\[14\] _03081_ _03398_ _03080_ VGND VGND VPWR VPWR _02428_ sky130_fd_sc_hd__o211a_1
X_11037_ net1872 _05683_ _06215_ VGND VGND VPWR VPWR _06222_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_108_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16894_ _04148_ per_uart.rx_avail _04138_ VGND VGND VPWR VPWR _04173_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_125_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15845_ _02757_ _03307_ _03316_ _03331_ _02846_ VGND VGND VPWR VPWR _03332_ sky130_fd_sc_hd__a311o_2
X_15776_ CPU.aluIn1\[10\] _02958_ _03241_ _03264_ _02995_ VGND VGND VPWR VPWR _02424_
+ sky130_fd_sc_hd__o221a_1
X_12988_ CPU.registerFile\[23\]\[3\] _07236_ _07239_ CPU.registerFile\[19\]\[3\] _07427_
+ VGND VGND VPWR VPWR _07428_ sky130_fd_sc_hd__o221a_1
XFILLER_0_148_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17515_ net704 _01803_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11939_ _06736_ VGND VGND VPWR VPWR _01601_ sky130_fd_sc_hd__clkbuf_1
X_17446_ net635 _01734_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13609_ CPU.registerFile\[31\]\[21\] _07772_ _07773_ CPU.registerFile\[27\]\[21\]
+ _08030_ VGND VGND VPWR VPWR _08031_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_41_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17377_ net566 _01665_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_888 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_131_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16328_ CPU.registerFile\[9\]\[27\] CPU.registerFile\[13\]\[27\] _02999_ VGND VGND
+ VPWR VPWR _03800_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16259_ CPU.registerFile\[8\]\[25\] _02894_ _02764_ _03732_ VGND VGND VPWR VPWR _03733_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_136_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09702_ _05391_ _04211_ _04219_ CPU.aluReg\[2\] _05392_ VGND VGND VPWR VPWR _05393_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_52_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09633_ _04918_ _05326_ VGND VGND VPWR VPWR _05327_ sky130_fd_sc_hd__or2_1
X_09564_ _04424_ _04405_ _04423_ VGND VGND VPWR VPWR _05260_ sky130_fd_sc_hd__nor3_1
X_08515_ CPU.rs2\[24\] _04201_ _04206_ VGND VGND VPWR VPWR _04235_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09495_ _04857_ _04890_ VGND VGND VPWR VPWR _05194_ sky130_fd_sc_hd__and2b_1
XFILLER_0_148_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_156_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10270_ _05516_ net2131 _05751_ VGND VGND VPWR VPWR _05754_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12911_ CPU.registerFile\[28\]\[1\] CPU.registerFile\[24\]\[1\] _07352_ VGND VGND
+ VPWR VPWR _07353_ sky130_fd_sc_hd__mux2_1
X_13891_ CPU.registerFile\[6\]\[30\] CPU.registerFile\[7\]\[30\] _07263_ VGND VGND
+ VPWR VPWR _08304_ sky130_fd_sc_hd__mux2_1
X_15190__103 clknet_1_1__leaf__02750_ VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__inv_2
X_15630_ CPU.registerFile\[15\]\[7\] CPU.registerFile\[11\]\[7\] _02773_ VGND VGND
+ VPWR VPWR _03122_ sky130_fd_sc_hd__mux2_1
X_12842_ _04971_ VGND VGND VPWR VPWR _07285_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_87_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_87_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _02797_ _03051_ _03052_ _03053_ _03054_ VGND VGND VPWR VPWR _03055_ sky130_fd_sc_hd__a221o_1
X_17300_ net489 _01588_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11724_ net4 _06574_ _06616_ _06607_ VGND VGND VPWR VPWR _01695_ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18280_ net113 _02560_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_25_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15492_ _05050_ _02986_ _02987_ VGND VGND VPWR VPWR _02988_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17231_ net421 _01519_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11655_ net1450 _06575_ _06578_ _06539_ VGND VGND VPWR VPWR _01726_ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17162_ net386 _01450_ VGND VGND VPWR VPWR CPU.aluReg\[26\] sky130_fd_sc_hd__dfxtp_1
X_10606_ mapped_spi_flash.rcv_data\[19\] _05981_ VGND VGND VPWR VPWR _05986_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14374_ clknet_1_0__leaf__02653_ VGND VGND VPWR VPWR _02654_ sky130_fd_sc_hd__buf_1
X_11586_ _06512_ _05923_ VGND VGND VPWR VPWR _06529_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16113_ _03015_ _03589_ _03590_ _03591_ _02930_ VGND VGND VPWR VPWR _03592_ sky130_fd_sc_hd__a221o_1
X_13325_ CPU.registerFile\[8\]\[12\] CPU.registerFile\[12\]\[12\] _07318_ VGND VGND
+ VPWR VPWR _07756_ sky130_fd_sc_hd__mux2_1
X_10537_ _05856_ _05937_ VGND VGND VPWR VPWR _05938_ sky130_fd_sc_hd__or2_1
X_17093_ net351 _01415_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_118_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__02751_ clknet_0__02751_ VGND VGND VPWR VPWR clknet_1_1__leaf__02751_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_134_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16044_ CPU.registerFile\[22\]\[18\] CPU.registerFile\[23\]\[18\] _03066_ VGND VGND
+ VPWR VPWR _03525_ sky130_fd_sc_hd__mux2_1
X_13256_ CPU.registerFile\[28\]\[10\] CPU.registerFile\[24\]\[10\] _07476_ VGND VGND
+ VPWR VPWR _07689_ sky130_fd_sc_hd__mux2_1
X_10468_ _04507_ _04551_ _04552_ VGND VGND VPWR VPWR _05880_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__02682_ clknet_0__02682_ VGND VGND VPWR VPWR clknet_1_1__leaf__02682_
+ sky130_fd_sc_hd__clkbuf_16
X_12207_ CPU.aluReg\[27\] CPU.aluReg\[25\] _06871_ VGND VGND VPWR VPWR _06889_ sky130_fd_sc_hd__mux2_1
X_13187_ CPU.registerFile\[15\]\[8\] _07325_ _07620_ _07621_ _07327_ VGND VGND VPWR
+ VPWR _07622_ sky130_fd_sc_hd__o221a_1
X_10399_ _05816_ _05828_ VGND VGND VPWR VPWR _05829_ sky130_fd_sc_hd__and2_1
X_12138_ _05188_ net1971 _06841_ VGND VGND VPWR VPWR _06842_ sky130_fd_sc_hd__mux2_1
X_17995_ clknet_leaf_10_clk _02279_ VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[9\]
+ sky130_fd_sc_hd__dfxtp_1
X_16946_ net241 _01272_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_12069_ _06782_ VGND VGND VPWR VPWR _06805_ sky130_fd_sc_hd__clkbuf_4
X_14567__684 clknet_1_1__leaf__02672_ VGND VGND VPWR VPWR net716 sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_1_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_8
X_16877_ per_uart.uart0.rx_count16\[2\] _04156_ per_uart.uart0.rx_count16\[3\] VGND
+ VGND VPWR VPWR _04161_ sky130_fd_sc_hd__a21o_1
X_15828_ _02885_ _03312_ _03313_ _03314_ _03054_ VGND VGND VPWR VPWR _03315_ sky130_fd_sc_hd__a221o_1
X_15002__1076 clknet_1_1__leaf__02715_ VGND VGND VPWR VPWR net1108 sky130_fd_sc_hd__inv_2
XFILLER_0_59_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15759_ CPU.registerFile\[15\]\[10\] CPU.registerFile\[11\]\[10\] _03247_ VGND VGND
+ VPWR VPWR _03248_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09280_ _04502_ VGND VGND VPWR VPWR _04989_ sky130_fd_sc_hd__buf_2
XFILLER_0_75_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17429_ net618 net1449 VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14732__832 clknet_1_1__leaf__02689_ VGND VGND VPWR VPWR net864 sky130_fd_sc_hd__inv_2
XFILLER_0_15_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_151_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload50 clknet_1_0__leaf__02711_ VGND VGND VPWR VPWR clkload50/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_140_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload61 clknet_1_1__leaf__02693_ VGND VGND VPWR VPWR clkload61/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload72 clknet_1_1__leaf__02674_ VGND VGND VPWR VPWR clkload72/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_3_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload83 clknet_1_0__leaf__02661_ VGND VGND VPWR VPWR clkload83/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload94 clknet_1_1__leaf__08465_ VGND VGND VPWR VPWR clkload94/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08995_ CPU.cycles\[29\] _04687_ _04712_ VGND VGND VPWR VPWR _04713_ sky130_fd_sc_hd__a21o_4
XTAP_TAPCELL_ROW_149_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09616_ mapped_spi_flash.rcv_data\[29\] _04709_ _05309_ VGND VGND VPWR VPWR _05310_
+ sky130_fd_sc_hd__a21o_1
X_09547_ _04273_ net1288 VGND VGND VPWR VPWR _05244_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09478_ CPU.cycles\[11\] _04989_ _04916_ _05177_ VGND VGND VPWR VPWR _05178_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_66_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14024__303 clknet_1_1__leaf__08362_ VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__inv_2
XFILLER_0_136_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14395__529 clknet_1_0__leaf__02655_ VGND VGND VPWR VPWR net561 sky130_fd_sc_hd__inv_2
XFILLER_0_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18373__32 VGND VGND VPWR VPWR _18373__32/HI net32 sky130_fd_sc_hd__conb_1
Xclkload0 clknet_2_0__leaf_clk VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__clkinv_2
X_11440_ _06436_ VGND VGND VPWR VPWR _01803_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11371_ _05495_ net2006 _06397_ VGND VGND VPWR VPWR _06400_ sky130_fd_sc_hd__mux2_1
X_13110_ _07232_ _07539_ _07546_ VGND VGND VPWR VPWR _07547_ sky130_fd_sc_hd__a21o_1
X_10322_ _05499_ net2072 _05777_ VGND VGND VPWR VPWR _05782_ sky130_fd_sc_hd__mux2_1
X_14090_ _04484_ net1273 VGND VGND VPWR VPWR _08371_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_885 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13041_ _04938_ VGND VGND VPWR VPWR _07480_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_30_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10253_ _05499_ net1941 _05740_ VGND VGND VPWR VPWR _05745_ sky130_fd_sc_hd__mux2_1
X_10184_ net2332 _05698_ _05692_ VGND VGND VPWR VPWR _05699_ sky130_fd_sc_hd__mux2_1
X_14861__949 clknet_1_1__leaf__02701_ VGND VGND VPWR VPWR net981 sky130_fd_sc_hd__inv_2
X_16800_ _04050_ _04107_ _04108_ _04109_ VGND VGND VPWR VPWR _04110_ sky130_fd_sc_hd__a31o_1
X_17780_ net969 _02064_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_89_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16731_ _04499_ VGND VGND VPWR VPWR _04052_ sky130_fd_sc_hd__clkbuf_2
X_13943_ net1479 _08018_ _08354_ _08017_ VGND VGND VPWR VPWR _01326_ sky130_fd_sc_hd__o211a_1
X_16662_ CPU.PC\[2\] _08379_ _08454_ VGND VGND VPWR VPWR _03993_ sky130_fd_sc_hd__or3b_1
X_13874_ _07260_ _08287_ VGND VGND VPWR VPWR _08288_ sky130_fd_sc_hd__or2_1
X_15613_ _02812_ _03102_ _03105_ _02948_ VGND VGND VPWR VPWR _03106_ sky130_fd_sc_hd__o211a_1
X_12825_ _04785_ VGND VGND VPWR VPWR _07268_ sky130_fd_sc_hd__buf_4
XFILLER_0_158_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18332_ clknet_leaf_6_clk _02612_ VGND VGND VPWR VPWR per_uart.uart0.tx_bitcount\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_15544_ CPU.registerFile\[12\]\[5\] _05049_ VGND VGND VPWR VPWR _03038_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11707_ mapped_spi_ram.rcv_data\[8\] _06601_ VGND VGND VPWR VPWR _06608_ sky130_fd_sc_hd__or2_1
X_18263_ clknet_leaf_2_clk _02543_ VGND VGND VPWR VPWR per_uart.uart0.rxd_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_15475_ _02858_ _02968_ _02970_ _02864_ VGND VGND VPWR VPWR _02971_ sky130_fd_sc_hd__a211o_1
X_12687_ CPU.cycles\[28\] CPU.cycles\[29\] _07170_ VGND VGND VPWR VPWR _07172_ sky130_fd_sc_hd__and3_1
X_17214_ net404 _01502_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18194_ net225 _02474_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_11638_ _06549_ _06564_ VGND VGND VPWR VPWR _06565_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17145_ net369 _01433_ VGND VGND VPWR VPWR CPU.aluReg\[9\] sky130_fd_sc_hd__dfxtp_1
X_11569_ _06493_ VGND VGND VPWR VPWR _06517_ sky130_fd_sc_hd__buf_2
XFILLER_0_123_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold707 CPU.registerFile\[26\]\[12\] VGND VGND VPWR VPWR net1948 sky130_fd_sc_hd__dlygate4sd3_1
Xhold718 CPU.registerFile\[12\]\[3\] VGND VGND VPWR VPWR net1959 sky130_fd_sc_hd__dlygate4sd3_1
X_13308_ _05338_ _07738_ VGND VGND VPWR VPWR _07739_ sky130_fd_sc_hd__or2_1
Xhold729 CPU.registerFile\[2\]\[17\] VGND VGND VPWR VPWR net1970 sky130_fd_sc_hd__dlygate4sd3_1
X_17076_ net334 _01398_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16027_ CPU.registerFile\[28\]\[18\] _03064_ VGND VGND VPWR VPWR _03508_ sky130_fd_sc_hd__or2_1
X_13239_ _07397_ _07665_ _07672_ _07424_ VGND VGND VPWR VPWR _07673_ sky130_fd_sc_hd__a31o_2
Xclkbuf_1_1__f__02665_ clknet_0__02665_ VGND VGND VPWR VPWR clknet_1_1__leaf__02665_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__02696_ _02696_ VGND VGND VPWR VPWR clknet_0__02696_ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_0__07223_ _07223_ VGND VGND VPWR VPWR clknet_0__07223_ sky130_fd_sc_hd__clkbuf_16
X_08780_ _04499_ VGND VGND VPWR VPWR _04500_ sky130_fd_sc_hd__inv_2
X_17978_ net1166 _02262_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[23\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_127_Right_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09401_ _04256_ _04683_ VGND VGND VPWR VPWR _05105_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09332_ _04445_ _04488_ _05038_ _04768_ VGND VGND VPWR VPWR _05039_ sky130_fd_sc_hd__a22o_1
XFILLER_0_158_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_80_Left_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09263_ _04782_ _04972_ net1277 VGND VGND VPWR VPWR _04973_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_157_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14320__461 clknet_1_1__leaf__08465_ VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__inv_2
X_09194_ _04828_ _04905_ VGND VGND VPWR VPWR _04906_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08978_ net1580 _04696_ _04668_ VGND VGND VPWR VPWR _04697_ sky130_fd_sc_hd__mux2_1
Xhold67 mapped_spi_ram.div_counter\[0\] VGND VGND VPWR VPWR net1308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 mapped_spi_ram.cmd_addr\[26\] VGND VGND VPWR VPWR net1319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 mapped_spi_ram.rcv_data\[5\] VGND VGND VPWR VPWR net1330 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10940_ _06170_ VGND VGND VPWR VPWR _02037_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__02754_ clknet_0__02754_ VGND VGND VPWR VPWR clknet_1_0__leaf__02754_
+ sky130_fd_sc_hd__clkbuf_16
X_12761__211 clknet_1_1__leaf__07224_ VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_67_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10871_ _06133_ VGND VGND VPWR VPWR _02069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_119_Left_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__02685_ clknet_0__02685_ VGND VGND VPWR VPWR clknet_1_0__leaf__02685_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12610_ net1513 net2 VGND VGND VPWR VPWR _07128_ sky130_fd_sc_hd__nand2_2
X_14403__536 clknet_1_0__leaf__02656_ VGND VGND VPWR VPWR net568 sky130_fd_sc_hd__inv_2
X_13590_ _07405_ _08009_ _08010_ _08012_ _07359_ VGND VGND VPWR VPWR _08013_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12541_ net1688 _04797_ _07085_ VGND VGND VPWR VPWR _07093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15260_ _02758_ VGND VGND VPWR VPWR _02759_ sky130_fd_sc_hd__buf_4
XFILLER_0_152_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12472_ _07056_ VGND VGND VPWR VPWR _01353_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11423_ _05547_ net1720 _06419_ VGND VGND VPWR VPWR _06427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_9 _02819_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14142_ _08404_ VGND VGND VPWR VPWR _08405_ sky130_fd_sc_hd__buf_4
X_11354_ _05547_ net2421 _06382_ VGND VGND VPWR VPWR _06390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15001__1075 clknet_1_1__leaf__02715_ VGND VGND VPWR VPWR net1107 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_128_Left_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10305_ _05551_ net1818 _05762_ VGND VGND VPWR VPWR _05772_ sky130_fd_sc_hd__mux2_1
X_11285_ _06353_ VGND VGND VPWR VPWR _01875_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_111_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10236_ net2179 _05733_ _05670_ VGND VGND VPWR VPWR _05734_ sky130_fd_sc_hd__mux2_1
X_13024_ CPU.registerFile\[3\]\[4\] _07373_ _07462_ _07376_ VGND VGND VPWR VPWR _07463_
+ sky130_fd_sc_hd__o211a_1
X_17901_ net1090 _02185_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[19\] sky130_fd_sc_hd__dfxtp_1
X_17832_ net1021 _02116_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_10167_ _04932_ VGND VGND VPWR VPWR _05687_ sky130_fd_sc_hd__buf_2
XFILLER_0_83_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17763_ net952 _02047_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10098_ _05646_ VGND VGND VPWR VPWR _02370_ sky130_fd_sc_hd__clkbuf_1
X_16714_ _04033_ _04037_ _05942_ VGND VGND VPWR VPWR _02589_ sky130_fd_sc_hd__o21a_1
XFILLER_0_107_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13926_ _08334_ _08337_ _07474_ VGND VGND VPWR VPWR _08338_ sky130_fd_sc_hd__a21oi_2
X_17694_ net883 _01982_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_137_Left_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16645_ clknet_1_1__leaf__07219_ VGND VGND VPWR VPWR _03989_ sky130_fd_sc_hd__buf_1
X_13857_ CPU.registerFile\[5\]\[29\] _07577_ _08270_ _07638_ VGND VGND VPWR VPWR _08271_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12808_ _07243_ _07248_ _07250_ VGND VGND VPWR VPWR _07251_ sky130_fd_sc_hd__mux2_2
X_14679__785 clknet_1_0__leaf__02683_ VGND VGND VPWR VPWR net817 sky130_fd_sc_hd__inv_2
X_13788_ CPU.rs2\[26\] _07705_ _08189_ _08204_ _07737_ VGND VGND VPWR VPWR _01321_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_123_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18315_ clknet_leaf_16_clk _02595_ VGND VGND VPWR VPWR CPU.PC\[15\] sky130_fd_sc_hd__dfxtp_2
X_15527_ _02806_ VGND VGND VPWR VPWR _03022_ sky130_fd_sc_hd__buf_4
X_14378__513 clknet_1_0__leaf__02654_ VGND VGND VPWR VPWR net545 sky130_fd_sc_hd__inv_2
XFILLER_0_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12739_ _07215_ net1713 _07205_ VGND VGND VPWR VPWR _07216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18246_ net87 _02526_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15458_ _02827_ _02953_ _02954_ VGND VGND VPWR VPWR _02955_ sky130_fd_sc_hd__o21a_1
XFILLER_0_72_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18177_ net208 _02457_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_15389_ _02777_ VGND VGND VPWR VPWR _02887_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_13_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold504 CPU.registerFile\[3\]\[18\] VGND VGND VPWR VPWR net1745 sky130_fd_sc_hd__dlygate4sd3_1
X_17128_ clknet_leaf_22_clk _00031_ VGND VGND VPWR VPWR CPU.cycles\[24\] sky130_fd_sc_hd__dfxtp_1
Xhold515 CPU.registerFile\[13\]\[26\] VGND VGND VPWR VPWR net1756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold526 CPU.registerFile\[22\]\[24\] VGND VGND VPWR VPWR net1767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 CPU.registerFile\[22\]\[16\] VGND VGND VPWR VPWR net1778 sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 CPU.registerFile\[29\]\[21\] VGND VGND VPWR VPWR net1789 sky130_fd_sc_hd__dlygate4sd3_1
X_09950_ _05505_ net1702 _05559_ VGND VGND VPWR VPWR _05567_ sky130_fd_sc_hd__mux2_1
X_17059_ net317 _01381_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[21\] sky130_fd_sc_hd__dfxtp_1
Xhold559 CPU.registerFile\[17\]\[31\] VGND VGND VPWR VPWR net1800 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__02717_ clknet_0__02717_ VGND VGND VPWR VPWR clknet_1_1__leaf__02717_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08901_ _04524_ net1272 VGND VGND VPWR VPWR _04621_ sky130_fd_sc_hd__xor2_4
Xclkbuf_0__02748_ _02748_ VGND VGND VPWR VPWR clknet_0__02748_ sky130_fd_sc_hd__clkbuf_16
X_09881_ _05089_ VGND VGND VPWR VPWR _05522_ sky130_fd_sc_hd__buf_4
X_14844__933 clknet_1_1__leaf__02700_ VGND VGND VPWR VPWR net965 sky130_fd_sc_hd__inv_2
XFILLER_0_148_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08832_ CPU.aluIn1\[13\] CPU.Bimm\[12\] VGND VGND VPWR VPWR _04552_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_0__02679_ _02679_ VGND VGND VPWR VPWR clknet_0__02679_ sky130_fd_sc_hd__clkbuf_16
Xhold1204 CPU.registerFile\[28\]\[25\] VGND VGND VPWR VPWR net2445 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_148_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1215 CPU.registerFile\[2\]\[7\] VGND VGND VPWR VPWR net2456 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1226 mapped_spi_flash.rcv_data\[12\] VGND VGND VPWR VPWR net2467 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1237 CPU.registerFile\[2\]\[8\] VGND VGND VPWR VPWR net2478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1248 CPU.registerFile\[11\]\[11\] VGND VGND VPWR VPWR net2489 sky130_fd_sc_hd__dlygate4sd3_1
X_08763_ CPU.Jimm\[14\] VGND VGND VPWR VPWR _04483_ sky130_fd_sc_hd__clkbuf_4
Xhold1259 CPU.registerFile\[8\]\[28\] VGND VGND VPWR VPWR net2500 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08694_ _04411_ _04300_ _04413_ VGND VGND VPWR VPWR _04414_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09315_ CPU.PC\[18\] _04926_ CPU.PC\[19\] VGND VGND VPWR VPWR _05023_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14890__975 clknet_1_1__leaf__02704_ VGND VGND VPWR VPWR net1007 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_62_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09246_ _04950_ _04941_ _04940_ _04956_ VGND VGND VPWR VPWR _04957_ sky130_fd_sc_hd__or4b_4
XTAP_TAPCELL_ROW_32_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09177_ CPU.PC\[9\] CPU.Bimm\[9\] _04820_ _04888_ VGND VGND VPWR VPWR _04889_ sky130_fd_sc_hd__a31o_1
XFILLER_0_133_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11070_ _06239_ VGND VGND VPWR VPWR _01976_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10021_ net1618 _04933_ _05596_ VGND VGND VPWR VPWR _05605_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11972_ _04780_ net1782 _06747_ VGND VGND VPWR VPWR _06754_ sky130_fd_sc_hd__mux2_1
X_13711_ CPU.registerFile\[8\]\[24\] CPU.registerFile\[12\]\[24\] _07339_ VGND VGND
+ VPWR VPWR _08130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10923_ _06161_ VGND VGND VPWR VPWR _02045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16430_ _03897_ _03898_ _02856_ VGND VGND VPWR VPWR _03899_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13642_ _08059_ _08062_ _07514_ VGND VGND VPWR VPWR _08063_ sky130_fd_sc_hd__a21oi_4
X_10854_ _06124_ VGND VGND VPWR VPWR _02077_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__02668_ clknet_0__02668_ VGND VGND VPWR VPWR clknet_1_0__leaf__02668_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16361_ CPU.registerFile\[8\]\[28\] _02789_ _02790_ _03831_ VGND VGND VPWR VPWR _03832_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13573_ CPU.registerFile\[16\]\[20\] CPU.registerFile\[20\]\[20\] _07648_ VGND VGND
+ VPWR VPWR _07996_ sky130_fd_sc_hd__mux2_1
X_10785_ _05524_ net1708 _06081_ VGND VGND VPWR VPWR _06088_ sky130_fd_sc_hd__mux2_1
X_18100_ net163 _02380_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15312_ _02795_ _02808_ _02810_ VGND VGND VPWR VPWR _02811_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_30_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12524_ _07083_ VGND VGND VPWR VPWR _01328_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16292_ CPU.registerFile\[8\]\[26\] CPU.registerFile\[12\]\[26\] _02798_ VGND VGND
+ VPWR VPWR _03765_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18031_ net1204 _02311_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12455_ _05448_ net2271 _07012_ VGND VGND VPWR VPWR _07047_ sky130_fd_sc_hd__mux2_1
X_15228__138 clknet_1_0__leaf__02753_ VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_97_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11406_ _05530_ net2081 _06408_ VGND VGND VPWR VPWR _06418_ sky130_fd_sc_hd__mux2_1
X_15174_ clknet_1_0__leaf__02720_ VGND VGND VPWR VPWR _02748_ sky130_fd_sc_hd__buf_1
XFILLER_0_1_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12386_ _07010_ VGND VGND VPWR VPWR _01393_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14002__283 clknet_1_0__leaf__08360_ VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__inv_2
X_14125_ _04782_ _05132_ _08387_ VGND VGND VPWR VPWR _08392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11337_ _05530_ net2343 _06371_ VGND VGND VPWR VPWR _06381_ sky130_fd_sc_hd__mux2_1
X_11268_ _06344_ VGND VGND VPWR VPWR _01883_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13007_ CPU.registerFile\[13\]\[3\] _07282_ _07446_ VGND VGND VPWR VPWR _07447_ sky130_fd_sc_hd__o21a_1
X_10219_ _05722_ VGND VGND VPWR VPWR _02325_ sky130_fd_sc_hd__clkbuf_1
X_11199_ _05528_ net1885 _06299_ VGND VGND VPWR VPWR _06308_ sky130_fd_sc_hd__mux2_1
X_17815_ net1004 _02099_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_128_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_145_Left_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17746_ net935 _02030_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[0\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13909_ _08317_ _08318_ _08319_ _08321_ _07359_ VGND VGND VPWR VPWR _08322_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_18_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17677_ net866 _01965_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16569__42 clknet_1_1__leaf__03968_ VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__inv_2
XFILLER_0_45_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09100_ _04497_ VGND VGND VPWR VPWR _04812_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_44_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16584__56 clknet_1_1__leaf__03969_ VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__inv_2
XFILLER_0_5_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_154_Left_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_878 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09031_ CPU.Bimm\[7\] _04498_ _04746_ VGND VGND VPWR VPWR _04747_ sky130_fd_sc_hd__a21o_2
XFILLER_0_150_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18229_ net70 _02509_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold301 CPU.aluShamt\[3\] VGND VGND VPWR VPWR net1542 sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 _04143_ VGND VGND VPWR VPWR net1553 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 CPU.registerFile\[5\]\[21\] VGND VGND VPWR VPWR net1564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 per_uart.uart0.txd_reg\[2\] VGND VGND VPWR VPWR net1575 sky130_fd_sc_hd__dlygate4sd3_1
Xhold345 CPU.registerFile\[6\]\[19\] VGND VGND VPWR VPWR net1586 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 per_uart.uart0.txd_reg\[4\] VGND VGND VPWR VPWR net1597 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 CPU.registerFile\[6\]\[29\] VGND VGND VPWR VPWR net1608 sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 CPU.registerFile\[12\]\[13\] VGND VGND VPWR VPWR net1619 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ _04661_ _04660_ VGND VGND VPWR VPWR _05557_ sky130_fd_sc_hd__nor2b_2
X_14432__562 clknet_1_1__leaf__02659_ VGND VGND VPWR VPWR net594 sky130_fd_sc_hd__inv_2
Xhold389 CPU.registerFile\[16\]\[2\] VGND VGND VPWR VPWR net1630 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09864_ _05510_ VGND VGND VPWR VPWR _02500_ sky130_fd_sc_hd__clkbuf_1
Xhold1001 CPU.registerFile\[19\]\[14\] VGND VGND VPWR VPWR net2242 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1012 CPU.registerFile\[23\]\[19\] VGND VGND VPWR VPWR net2253 sky130_fd_sc_hd__dlygate4sd3_1
X_08815_ _04522_ _04534_ _04520_ _04517_ CPU.aluIn1\[4\] VGND VGND VPWR VPWR _04535_
+ sky130_fd_sc_hd__a32o_1
Xhold1023 CPU.registerFile\[8\]\[22\] VGND VGND VPWR VPWR net2264 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1034 CPU.registerFile\[28\]\[28\] VGND VGND VPWR VPWR net2275 sky130_fd_sc_hd__dlygate4sd3_1
X_09795_ _05468_ VGND VGND VPWR VPWR _02527_ sky130_fd_sc_hd__clkbuf_1
Xhold1045 CPU.registerFile\[2\]\[16\] VGND VGND VPWR VPWR net2286 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1056 CPU.registerFile\[6\]\[17\] VGND VGND VPWR VPWR net2297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 CPU.registerFile\[13\]\[11\] VGND VGND VPWR VPWR net2308 sky130_fd_sc_hd__dlygate4sd3_1
X_08746_ _04356_ VGND VGND VPWR VPWR _04466_ sky130_fd_sc_hd__inv_2
Xhold1078 CPU.registerFile\[8\]\[7\] VGND VGND VPWR VPWR net2319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1089 mapped_spi_flash.rcv_data\[15\] VGND VGND VPWR VPWR net2330 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_207 _07914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_218 clknet_2_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08677_ CPU.aluIn1\[12\] VGND VGND VPWR VPWR _04397_ sky130_fd_sc_hd__inv_2
XANTENNA_229 clknet_1_1__leaf__02693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15000__1074 clknet_1_1__leaf__02715_ VGND VGND VPWR VPWR net1106 sky130_fd_sc_hd__inv_2
XFILLER_0_138_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_875 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10570_ net1551 mapped_spi_flash.state\[3\] VGND VGND VPWR VPWR _05962_ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09229_ _04782_ _04939_ net1277 VGND VGND VPWR VPWR _04940_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12240_ CPU.aluReg\[19\] _06914_ _06891_ VGND VGND VPWR VPWR _06915_ sky130_fd_sc_hd__mux2_1
X_14515__637 clknet_1_0__leaf__02667_ VGND VGND VPWR VPWR net669 sky130_fd_sc_hd__inv_2
X_12171_ _06855_ _06857_ _06862_ VGND VGND VPWR VPWR _01494_ sky130_fd_sc_hd__o21a_1
XFILLER_0_20_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14253__425 clknet_1_0__leaf__08435_ VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__inv_2
X_11122_ _06267_ VGND VGND VPWR VPWR _01952_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_92_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold890 CPU.registerFile\[20\]\[19\] VGND VGND VPWR VPWR net2131 sky130_fd_sc_hd__dlygate4sd3_1
X_11053_ _06230_ VGND VGND VPWR VPWR _01984_ sky130_fd_sc_hd__clkbuf_1
X_15930_ CPU.registerFile\[28\]\[15\] CPU.registerFile\[24\]\[15\] _02881_ VGND VGND
+ VPWR VPWR _03414_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10004_ _05595_ VGND VGND VPWR VPWR _05596_ sky130_fd_sc_hd__buf_4
X_15861_ CPU.registerFile\[29\]\[13\] _02800_ VGND VGND VPWR VPWR _03347_ sky130_fd_sc_hd__or2_1
X_17600_ net789 _01888_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_15792_ _02777_ VGND VGND VPWR VPWR _03280_ sky130_fd_sc_hd__buf_4
X_17531_ net720 _01819_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_11955_ _06744_ VGND VGND VPWR VPWR _01593_ sky130_fd_sc_hd__clkbuf_1
X_14561__679 clknet_1_0__leaf__02671_ VGND VGND VPWR VPWR net711 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_123_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10906_ _06152_ VGND VGND VPWR VPWR _02053_ sky130_fd_sc_hd__clkbuf_1
X_17462_ net651 _01750_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11886_ CPU.registerFile\[10\]\[1\] _05733_ _06674_ VGND VGND VPWR VPWR _06708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16413_ CPU.registerFile\[9\]\[29\] _08404_ _02860_ VGND VGND VPWR VPWR _03883_ sky130_fd_sc_hd__o21a_1
X_13625_ _07379_ _08042_ _08046_ _07268_ VGND VGND VPWR VPWR _08047_ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10837_ _06115_ VGND VGND VPWR VPWR _02085_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17393_ net582 _01681_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[25\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16344_ CPU.registerFile\[17\]\[27\] CPU.registerFile\[21\]\[27\] _05405_ VGND VGND
+ VPWR VPWR _03816_ sky130_fd_sc_hd__mux2_1
X_13556_ CPU.registerFile\[30\]\[19\] CPU.registerFile\[26\]\[19\] _04937_ VGND VGND
+ VPWR VPWR _07980_ sky130_fd_sc_hd__mux2_1
X_10768_ _05507_ net1596 _06070_ VGND VGND VPWR VPWR _06079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12507_ net1905 _05719_ _07071_ VGND VGND VPWR VPWR _07075_ sky130_fd_sc_hd__mux2_1
X_16275_ CPU.registerFile\[19\]\[25\] _05071_ _02873_ _03748_ VGND VGND VPWR VPWR
+ _03749_ sky130_fd_sc_hd__o211a_1
X_13487_ _07351_ _07912_ VGND VGND VPWR VPWR _07913_ sky130_fd_sc_hd__or2_1
X_10699_ _06042_ VGND VGND VPWR VPWR _02150_ sky130_fd_sc_hd__clkbuf_1
X_18014_ net1187 _02294_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_12438_ _07038_ VGND VGND VPWR VPWR _01369_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_669 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12369_ _05230_ net2434 _06999_ VGND VGND VPWR VPWR _07002_ sky130_fd_sc_hd__mux2_1
X_14108_ _08382_ VGND VGND VPWR VPWR _01463_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15088_ net1423 _07182_ VGND VGND VPWR VPWR _02731_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08600_ CPU.rs2\[11\] _04199_ _04204_ VGND VGND VPWR VPWR _04320_ sky130_fd_sc_hd__a21o_1
X_09580_ _04484_ _04624_ VGND VGND VPWR VPWR _05275_ sky130_fd_sc_hd__or2_2
XFILLER_0_54_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08531_ CPU.rs2\[17\] _04200_ _04205_ VGND VGND VPWR VPWR _04251_ sky130_fd_sc_hd__a21oi_1
X_17729_ net918 _02013_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_46_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_154_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_154_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09014_ _04730_ VGND VGND VPWR VPWR _04731_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold120 mapped_spi_ram.cmd_addr\[16\] VGND VGND VPWR VPWR net1361 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 mapped_spi_ram.cmd_addr\[10\] VGND VGND VPWR VPWR net1372 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 mapped_spi_flash.cmd_addr\[10\] VGND VGND VPWR VPWR net1383 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold153 mapped_spi_ram.cmd_addr\[21\] VGND VGND VPWR VPWR net1394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 _02192_ VGND VGND VPWR VPWR net1405 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold175 CPU.cycles\[17\] VGND VGND VPWR VPWR net1416 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold186 _00039_ VGND VGND VPWR VPWR net1427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 _07165_ VGND VGND VPWR VPWR net1438 sky130_fd_sc_hd__dlygate4sd3_1
X_09916_ _05545_ net2515 _05533_ VGND VGND VPWR VPWR _05546_ sky130_fd_sc_hd__mux2_1
X_09847_ _04747_ VGND VGND VPWR VPWR _05499_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14703__807 clknet_1_0__leaf__02685_ VGND VGND VPWR VPWR net839 sky130_fd_sc_hd__inv_2
X_15257__164 clknet_1_1__leaf__02756_ VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__inv_2
X_09778_ _05459_ VGND VGND VPWR VPWR _02535_ sky130_fd_sc_hd__clkbuf_1
X_08729_ _04446_ _04387_ _04448_ VGND VGND VPWR VPWR _04449_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_1_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ mapped_spi_ram.rcv_bitcount\[4\] _06571_ VGND VGND VPWR VPWR _06629_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_789 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16548__23 clknet_1_0__leaf__03966_ VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__inv_2
X_11671_ mapped_spi_ram.rcv_data\[23\] _06577_ VGND VGND VPWR VPWR _06587_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13410_ CPU.registerFile\[16\]\[15\] CPU.registerFile\[20\]\[15\] _07233_ VGND VGND
+ VPWR VPWR _07838_ sky130_fd_sc_hd__mux2_1
X_10622_ mapped_spi_flash.rcv_data\[12\] _05994_ VGND VGND VPWR VPWR _05995_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13341_ CPU.registerFile\[15\]\[13\] _07629_ _07488_ CPU.registerFile\[11\]\[13\]
+ _07770_ VGND VGND VPWR VPWR _07771_ sky130_fd_sc_hd__o221a_1
XFILLER_0_64_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16563__37 clknet_1_0__leaf__03967_ VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__inv_2
XFILLER_0_134_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10553_ _05948_ net2338 _05950_ VGND VGND VPWR VPWR _05951_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16060_ _03022_ _03537_ _03538_ _03539_ _03028_ VGND VGND VPWR VPWR _03540_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_20_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13272_ net2428 _07358_ _07688_ _07704_ _05844_ VGND VGND VPWR VPWR _01305_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_94_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10484_ _04548_ _05893_ VGND VGND VPWR VPWR _05894_ sky130_fd_sc_hd__xnor2_1
X_12223_ CPU.aluReg\[23\] _06901_ _06891_ VGND VGND VPWR VPWR _06902_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12154_ _05381_ net2304 _06841_ VGND VGND VPWR VPWR _06850_ sky130_fd_sc_hd__mux2_1
X_11105_ _06258_ VGND VGND VPWR VPWR _01960_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_9_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16962_ net257 _01288_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_12085_ _06813_ VGND VGND VPWR VPWR _01531_ sky130_fd_sc_hd__clkbuf_1
X_11036_ _06221_ VGND VGND VPWR VPWR _01992_ sky130_fd_sc_hd__clkbuf_1
X_15913_ _08407_ _03374_ _03383_ _03397_ _02846_ VGND VGND VPWR VPWR _03398_ sky130_fd_sc_hd__a311o_2
X_16893_ _04171_ _04170_ _04172_ _03632_ VGND VGND VPWR VPWR _02633_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_108_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15844_ _02936_ _03323_ _03330_ _02934_ VGND VGND VPWR VPWR _03331_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15775_ _08408_ _03253_ _03263_ _02993_ VGND VGND VPWR VPWR _03264_ sky130_fd_sc_hd__a31o_1
X_12987_ _05338_ _07426_ VGND VGND VPWR VPWR _07427_ sky130_fd_sc_hd__or2_1
X_17514_ net703 _01802_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_11938_ CPU.registerFile\[11\]\[9\] _05717_ _06733_ VGND VGND VPWR VPWR _06736_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_918 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17445_ net634 _01733_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11869_ _06699_ VGND VGND VPWR VPWR _01634_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13608_ _07370_ _08029_ VGND VGND VPWR VPWR _08030_ sky130_fd_sc_hd__or2_1
X_17376_ net565 _01664_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_41_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_227 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16327_ _03015_ _03796_ _03797_ _03798_ _08396_ VGND VGND VPWR VPWR _03799_ sky130_fd_sc_hd__a221o_1
X_13539_ CPU.registerFile\[1\]\[19\] _07576_ _07962_ _07639_ VGND VGND VPWR VPWR _07963_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16258_ CPU.registerFile\[12\]\[25\] _05049_ VGND VGND VPWR VPWR _03732_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16189_ CPU.aluIn1\[22\] _02958_ _03650_ _03665_ _02995_ VGND VGND VPWR VPWR _02436_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09701_ _04306_ _04683_ VGND VGND VPWR VPWR _05392_ sky130_fd_sc_hd__nor2_1
X_14979__1055 clknet_1_1__leaf__02713_ VGND VGND VPWR VPWR net1087 sky130_fd_sc_hd__inv_2
XFILLER_0_156_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09632_ CPU.PC\[5\] _04917_ VGND VGND VPWR VPWR _05326_ sky130_fd_sc_hd__nor2_1
XFILLER_0_156_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14544__663 clknet_1_0__leaf__02670_ VGND VGND VPWR VPWR net695 sky130_fd_sc_hd__inv_2
X_09563_ _04919_ _05258_ VGND VGND VPWR VPWR _05259_ sky130_fd_sc_hd__or2_1
X_08514_ CPU.aluIn1\[25\] _04233_ VGND VGND VPWR VPWR _04234_ sky130_fd_sc_hd__nand2_1
X_09494_ _04716_ _05192_ _04717_ VGND VGND VPWR VPWR _05193_ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_156_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14627__738 clknet_1_1__leaf__02678_ VGND VGND VPWR VPWR net770 sky130_fd_sc_hd__inv_2
X_12910_ _04937_ VGND VGND VPWR VPWR _07352_ sky130_fd_sc_hd__clkbuf_8
X_13890_ CPU.registerFile\[2\]\[30\] CPU.registerFile\[3\]\[30\] _07263_ VGND VGND
+ VPWR VPWR _08303_ sky130_fd_sc_hd__mux2_1
X_12841_ CPU.registerFile\[8\]\[0\] CPU.registerFile\[12\]\[0\] _05284_ VGND VGND
+ VPWR VPWR _07284_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_100_Left_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15560_ _02806_ VGND VGND VPWR VPWR _03054_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_103_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11723_ mapped_spi_ram.rcv_data\[0\] _06576_ VGND VGND VPWR VPWR _06616_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15491_ CPU.registerFile\[16\]\[3\] _02832_ _02835_ CPU.registerFile\[17\]\[3\] _02940_
+ VGND VGND VPWR VPWR _02987_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_25_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ net420 _01518_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11654_ mapped_spi_ram.rcv_data\[31\] _06577_ VGND VGND VPWR VPWR _06578_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17161_ net385 _01449_ VGND VGND VPWR VPWR CPU.aluReg\[25\] sky130_fd_sc_hd__dfxtp_1
X_10605_ net2095 _05983_ _05985_ _05980_ VGND VGND VPWR VPWR _02186_ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14373_ clknet_1_0__leaf__07222_ VGND VGND VPWR VPWR _02653_ sky130_fd_sc_hd__buf_1
X_11585_ net1378 _06524_ _06528_ _06516_ VGND VGND VPWR VPWR _01746_ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16112_ CPU.registerFile\[27\]\[20\] _02928_ _02923_ VGND VGND VPWR VPWR _03591_
+ sky130_fd_sc_hd__o21a_1
X_13324_ _07273_ _07753_ _07754_ VGND VGND VPWR VPWR _07755_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17092_ net350 _01414_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[22\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__02750_ clknet_0__02750_ VGND VGND VPWR VPWR clknet_1_1__leaf__02750_
+ sky130_fd_sc_hd__clkbuf_16
X_10536_ mapped_spi_flash.cmd_addr\[1\] _04639_ _05820_ VGND VGND VPWR VPWR _05937_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16043_ _03065_ _03522_ _03523_ VGND VGND VPWR VPWR _03524_ sky130_fd_sc_hd__o21a_1
X_13255_ _07680_ _07687_ _07395_ VGND VGND VPWR VPWR _07688_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_108_Right_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__02681_ clknet_0__02681_ VGND VGND VPWR VPWR clknet_1_1__leaf__02681_
+ sky130_fd_sc_hd__clkbuf_16
X_10467_ net1368 _05849_ _05879_ _05855_ VGND VGND VPWR VPWR _02218_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12206_ _06888_ VGND VGND VPWR VPWR _01451_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13186_ _07311_ VGND VGND VPWR VPWR _07621_ sky130_fd_sc_hd__buf_4
X_10398_ mapped_spi_flash.cmd_addr\[30\] _05825_ _05827_ net11 VGND VGND VPWR VPWR
+ _05828_ sky130_fd_sc_hd__a22o_1
X_12137_ _06818_ VGND VGND VPWR VPWR _06841_ sky130_fd_sc_hd__clkbuf_4
X_17994_ clknet_leaf_10_clk _02278_ VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16945_ net240 _01271_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_12068_ _06804_ VGND VGND VPWR VPWR _01539_ sky130_fd_sc_hd__clkbuf_1
X_11019_ net1555 _05733_ _06178_ VGND VGND VPWR VPWR _06212_ sky130_fd_sc_hd__mux2_1
X_16876_ _04158_ _04160_ _05815_ VGND VGND VPWR VPWR _02628_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15827_ CPU.registerFile\[25\]\[12\] _03280_ _02803_ VGND VGND VPWR VPWR _03314_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_150_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15758_ _02760_ VGND VGND VPWR VPWR _03247_ sky130_fd_sc_hd__buf_4
XFILLER_0_129_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15689_ CPU.registerFile\[2\]\[8\] _02821_ _02813_ CPU.registerFile\[3\]\[8\] _05070_
+ VGND VGND VPWR VPWR _03180_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_390 _07285_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17428_ net617 _01716_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[21\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_138_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17359_ net548 _01647_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[23\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_151_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16542__18 clknet_1_0__leaf__03965_ VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__inv_2
XFILLER_0_42_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload40 clknet_1_0__leaf__02745_ VGND VGND VPWR VPWR clkload40/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_141_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload51 clknet_1_1__leaf__02710_ VGND VGND VPWR VPWR clkload51/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload62 clknet_1_1__leaf__02692_ VGND VGND VPWR VPWR clkload62/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_11_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload73 clknet_1_1__leaf__02673_ VGND VGND VPWR VPWR clkload73/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_140_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload84 clknet_1_1__leaf__02660_ VGND VGND VPWR VPWR clkload84/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_141_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload95 clknet_1_0__leaf__08464_ VGND VGND VPWR VPWR clkload95/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_3_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08994_ CPU.Bimm\[9\] _04498_ _04708_ _04707_ _04711_ VGND VGND VPWR VPWR _04712_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_149_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09615_ mapped_spi_ram.rcv_data\[29\] net17 _04643_ per_uart.rx_data\[5\] VGND VGND
+ VPWR VPWR _05309_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09546_ _04271_ _04211_ _04219_ CPU.aluReg\[8\] _05242_ VGND VGND VPWR VPWR _05243_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09477_ _04922_ _05176_ VGND VGND VPWR VPWR _05177_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14815__908 clknet_1_0__leaf__02696_ VGND VGND VPWR VPWR net940 sky130_fd_sc_hd__inv_2
X_14208__385 clknet_1_1__leaf__08430_ VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_22_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload1 clknet_2_2__leaf_clk VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_34_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12755__208 clknet_1_1__leaf__07221_ VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__inv_2
XFILLER_0_117_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11370_ _06399_ VGND VGND VPWR VPWR _01836_ sky130_fd_sc_hd__clkbuf_1
X_10321_ _05781_ VGND VGND VPWR VPWR _02267_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13040_ _07475_ _07477_ _07478_ VGND VGND VPWR VPWR _07479_ sky130_fd_sc_hd__o21a_1
X_10252_ _05744_ VGND VGND VPWR VPWR _02314_ sky130_fd_sc_hd__clkbuf_1
X_10183_ _05045_ VGND VGND VPWR VPWR _05698_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13942_ _07394_ _08339_ _08353_ _08015_ VGND VGND VPWR VPWR _08354_ sky130_fd_sc_hd__a211o_1
X_16730_ _04027_ _04039_ _05166_ VGND VGND VPWR VPWR _04051_ sky130_fd_sc_hd__a21o_1
X_16661_ _03991_ net2115 VGND VGND VPWR VPWR _03992_ sky130_fd_sc_hd__nand2_1
X_13873_ CPU.registerFile\[30\]\[29\] CPU.registerFile\[26\]\[29\] _07292_ VGND VGND
+ VPWR VPWR _08287_ sky130_fd_sc_hd__mux2_1
X_15612_ _02818_ _03103_ _03104_ VGND VGND VPWR VPWR _03105_ sky130_fd_sc_hd__a21o_1
X_12824_ _04939_ _07261_ _07266_ _04972_ VGND VGND VPWR VPWR _07267_ sky130_fd_sc_hd__a211o_1
XFILLER_0_69_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18331_ clknet_leaf_6_clk _02611_ VGND VGND VPWR VPWR per_uart.uart0.tx_bitcount\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15543_ CPU.registerFile\[14\]\[5\] CPU.registerFile\[10\]\[5\] _02761_ VGND VGND
+ VPWR VPWR _03037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11706_ net2485 _06603_ _06606_ _06607_ VGND VGND VPWR VPWR _01704_ sky130_fd_sc_hd__o211a_1
X_18262_ clknet_leaf_2_clk _02542_ VGND VGND VPWR VPWR per_uart.uart0.rxd_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_15474_ CPU.registerFile\[24\]\[3\] _02816_ _05071_ _02969_ VGND VGND VPWR VPWR _02970_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12686_ net1510 _07170_ VGND VGND VPWR VPWR _00035_ sky130_fd_sc_hd__xor2_1
XFILLER_0_53_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17213_ net403 _01501_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_14978__1054 clknet_1_0__leaf__02713_ VGND VGND VPWR VPWR net1086 sky130_fd_sc_hd__inv_2
X_18193_ net224 _02473_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_11637_ mapped_spi_ram.snd_bitcount\[1\] mapped_spi_ram.snd_bitcount\[0\] mapped_spi_ram.snd_bitcount\[2\]
+ VGND VGND VPWR VPWR _06564_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17144_ net368 _01432_ VGND VGND VPWR VPWR CPU.aluReg\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_499 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11568_ net1370 _06495_ _06514_ _06516_ VGND VGND VPWR VPWR _01751_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_133_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold708 CPU.registerFile\[24\]\[13\] VGND VGND VPWR VPWR net1949 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_133_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13307_ CPU.registerFile\[18\]\[12\] CPU.registerFile\[22\]\[12\] _07240_ VGND VGND
+ VPWR VPWR _07738_ sky130_fd_sc_hd__mux2_1
X_17075_ net333 _01397_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_10519_ _05886_ _05923_ VGND VGND VPWR VPWR _05924_ sky130_fd_sc_hd__nor2_1
Xhold719 CPU.registerFile\[23\]\[2\] VGND VGND VPWR VPWR net1960 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11499_ _05555_ net2102 _06432_ VGND VGND VPWR VPWR _06467_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16026_ CPU.registerFile\[30\]\[18\] CPU.registerFile\[26\]\[18\] _03247_ VGND VGND
+ VPWR VPWR _03507_ sky130_fd_sc_hd__mux2_1
X_13238_ _07411_ _07668_ _07671_ VGND VGND VPWR VPWR _07672_ sky130_fd_sc_hd__or3_1
Xclkbuf_1_1__f__02664_ clknet_0__02664_ VGND VGND VPWR VPWR clknet_1_1__leaf__02664_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_21_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__02695_ _02695_ VGND VGND VPWR VPWR clknet_0__02695_ sky130_fd_sc_hd__clkbuf_16
X_13169_ CPU.registerFile\[23\]\[8\] _07362_ _07363_ CPU.registerFile\[19\]\[8\] _07603_
+ VGND VGND VPWR VPWR _07604_ sky130_fd_sc_hd__o221a_1
Xclkbuf_0__07222_ _07222_ VGND VGND VPWR VPWR clknet_0__07222_ sky130_fd_sc_hd__clkbuf_16
X_17977_ net1165 _02261_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16859_ net1519 VGND VGND VPWR VPWR _04148_ sky130_fd_sc_hd__inv_2
X_09400_ _04439_ _04806_ VGND VGND VPWR VPWR _05104_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09331_ _05035_ _05037_ _04373_ VGND VGND VPWR VPWR _05038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09262_ _04971_ VGND VGND VPWR VPWR _04972_ sky130_fd_sc_hd__buf_6
XFILLER_0_117_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14656__764 clknet_1_1__leaf__02681_ VGND VGND VPWR VPWR net796 sky130_fd_sc_hd__inv_2
XFILLER_0_145_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09193_ _04835_ _04904_ _04833_ VGND VGND VPWR VPWR _04905_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_105_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08977_ _04695_ VGND VGND VPWR VPWR _04696_ sky130_fd_sc_hd__clkbuf_4
X_14821__912 clknet_1_0__leaf__02698_ VGND VGND VPWR VPWR net944 sky130_fd_sc_hd__inv_2
Xhold68 _06618_ VGND VGND VPWR VPWR net1309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 mapped_spi_flash.rcv_bitcount\[5\] VGND VGND VPWR VPWR net1320 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__02753_ clknet_0__02753_ VGND VGND VPWR VPWR clknet_1_0__leaf__02753_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_67_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10870_ net2456 _05721_ _06128_ VGND VGND VPWR VPWR _06133_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_84_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__02684_ clknet_0__02684_ VGND VGND VPWR VPWR clknet_1_0__leaf__02684_
+ sky130_fd_sc_hd__clkbuf_16
X_14739__839 clknet_1_0__leaf__02689_ VGND VGND VPWR VPWR net871 sky130_fd_sc_hd__inv_2
X_09529_ CPU.cycles\[9\] _04989_ VGND VGND VPWR VPWR _05227_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12540_ _07092_ VGND VGND VPWR VPWR _01288_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12471_ net1925 _05683_ _07049_ VGND VGND VPWR VPWR _07056_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11422_ _06426_ VGND VGND VPWR VPWR _01811_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14141_ _08403_ VGND VGND VPWR VPWR _08404_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_115_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11353_ _06389_ VGND VGND VPWR VPWR _01843_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10304_ _05771_ VGND VGND VPWR VPWR _02289_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11284_ CPU.registerFile\[9\]\[5\] _05725_ _06346_ VGND VGND VPWR VPWR _06353_ sky130_fd_sc_hd__mux2_1
X_13023_ CPU.registerFile\[2\]\[4\] _07374_ VGND VGND VPWR VPWR _07462_ sky130_fd_sc_hd__or2_1
X_17900_ net1089 _02184_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[18\] sky130_fd_sc_hd__dfxtp_1
X_10235_ _05425_ VGND VGND VPWR VPWR _05733_ sky130_fd_sc_hd__buf_2
X_17831_ net1020 _02115_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_10166_ _05686_ VGND VGND VPWR VPWR _02342_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17762_ net951 _02046_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_10097_ net1695 _05008_ _05644_ VGND VGND VPWR VPWR _05646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16713_ _04001_ _04034_ _04035_ _04036_ _07123_ VGND VGND VPWR VPWR _04037_ sky130_fd_sc_hd__o311a_1
X_13925_ _07650_ _08335_ _08336_ VGND VGND VPWR VPWR _08337_ sky130_fd_sc_hd__o21ai_1
X_17693_ net882 _01981_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13856_ CPU.registerFile\[4\]\[29\] _07374_ VGND VGND VPWR VPWR _08270_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12807_ _07249_ VGND VGND VPWR VPWR _07250_ sky130_fd_sc_hd__clkbuf_8
X_13787_ _07306_ _08196_ _08203_ _07703_ VGND VGND VPWR VPWR _08204_ sky130_fd_sc_hd__a31o_1
X_10999_ net2013 _05712_ _06201_ VGND VGND VPWR VPWR _06202_ sky130_fd_sc_hd__mux2_1
X_18314_ clknet_leaf_16_clk _02594_ VGND VGND VPWR VPWR CPU.PC\[14\] sky130_fd_sc_hd__dfxtp_2
X_15526_ _02848_ _03014_ _03020_ _02843_ VGND VGND VPWR VPWR _03021_ sky130_fd_sc_hd__a211o_1
X_12738_ per_uart.d_in_uart\[1\] _07178_ _07203_ per_uart.uart0.txd_reg\[2\] VGND
+ VGND VPWR VPWR _07215_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18245_ net86 _02525_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_15457_ CPU.registerFile\[18\]\[2\] _02832_ _02835_ CPU.registerFile\[19\]\[2\] _02796_
+ VGND VGND VPWR VPWR _02954_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_13_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12669_ CPU.cycles\[21\] _07160_ VGND VGND VPWR VPWR _07162_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_902 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18176_ net207 _02456_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_15388_ CPU.registerFile\[25\]\[1\] CPU.registerFile\[29\]\[1\] _02798_ VGND VGND
+ VPWR VPWR _02886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17127_ clknet_leaf_17_clk _00030_ VGND VGND VPWR VPWR CPU.cycles\[23\] sky130_fd_sc_hd__dfxtp_1
Xhold505 CPU.registerFile\[30\]\[6\] VGND VGND VPWR VPWR net1746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold516 CPU.registerFile\[20\]\[21\] VGND VGND VPWR VPWR net1757 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold527 per_uart.d_in_uart\[0\] VGND VGND VPWR VPWR net1768 sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 CPU.registerFile\[26\]\[16\] VGND VGND VPWR VPWR net1779 sky130_fd_sc_hd__dlygate4sd3_1
X_15205__117 clknet_1_0__leaf__02751_ VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__inv_2
X_17058_ net316 _01380_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[20\] sky130_fd_sc_hd__dfxtp_1
Xhold549 CPU.registerFile\[13\]\[0\] VGND VGND VPWR VPWR net1790 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__02716_ clknet_0__02716_ VGND VGND VPWR VPWR clknet_1_1__leaf__02716_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16009_ _03015_ _03488_ _03489_ _03490_ _02930_ VGND VGND VPWR VPWR _03491_ sky130_fd_sc_hd__a221o_1
XFILLER_0_110_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08900_ mapped_spi_ram.rcv_data\[23\] _04614_ _04618_ mapped_spi_flash.rcv_data\[23\]
+ VGND VGND VPWR VPWR _04620_ sky130_fd_sc_hd__a22oi_4
Xclkbuf_0__02747_ _02747_ VGND VGND VPWR VPWR clknet_0__02747_ sky130_fd_sc_hd__clkbuf_16
X_09880_ _05521_ VGND VGND VPWR VPWR _02495_ sky130_fd_sc_hd__clkbuf_1
X_08831_ _04550_ _04509_ VGND VGND VPWR VPWR _04551_ sky130_fd_sc_hd__or2_4
XFILLER_0_148_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__02678_ _02678_ VGND VGND VPWR VPWR clknet_0__02678_ sky130_fd_sc_hd__clkbuf_16
Xhold1205 CPU.registerFile\[22\]\[9\] VGND VGND VPWR VPWR net2446 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1216 CPU.registerFile\[31\]\[29\] VGND VGND VPWR VPWR net2457 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _04478_ _04480_ _04370_ VGND VGND VPWR VPWR _04482_ sky130_fd_sc_hd__o21ai_1
Xhold1227 CPU.registerFile\[24\]\[9\] VGND VGND VPWR VPWR net2468 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1238 CPU.aluReg\[28\] VGND VGND VPWR VPWR net2479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1249 mapped_spi_ram.rcv_data\[14\] VGND VGND VPWR VPWR net2490 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08693_ CPU.mem_wdata\[0\] _04203_ _04301_ _04412_ VGND VGND VPWR VPWR _04413_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15251__159 clknet_1_1__leaf__02755_ VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__inv_2
XFILLER_0_138_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09314_ _04835_ _04904_ VGND VGND VPWR VPWR _05022_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_158_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09245_ _04818_ _04952_ _04954_ _04955_ VGND VGND VPWR VPWR _04956_ sky130_fd_sc_hd__o22a_1
XFILLER_0_91_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09176_ _04859_ _04887_ VGND VGND VPWR VPWR _04888_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10020_ _05604_ VGND VGND VPWR VPWR _02406_ sky130_fd_sc_hd__clkbuf_1
X_14977__1053 clknet_1_0__leaf__02713_ VGND VGND VPWR VPWR net1085 sky130_fd_sc_hd__inv_2
XFILLER_0_98_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11971_ _06753_ VGND VGND VPWR VPWR _01586_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13710_ _07818_ _08127_ _08128_ VGND VGND VPWR VPWR _08129_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10922_ net1576 _05704_ _06154_ VGND VGND VPWR VPWR _06161_ sky130_fd_sc_hd__mux2_1
X_14327__468 clknet_1_0__leaf__08465_ VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__inv_2
X_13641_ _07650_ _08060_ _08061_ VGND VGND VPWR VPWR _08062_ sky130_fd_sc_hd__o21ai_1
X_10853_ net1847 _05704_ _06117_ VGND VGND VPWR VPWR _06124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__02667_ clknet_0__02667_ VGND VGND VPWR VPWR clknet_1_0__leaf__02667_
+ sky130_fd_sc_hd__clkbuf_16
X_16360_ CPU.registerFile\[12\]\[28\] _02791_ VGND VGND VPWR VPWR _03831_ sky130_fd_sc_hd__or2_1
X_13572_ CPU.registerFile\[23\]\[20\] _07282_ _07994_ VGND VGND VPWR VPWR _07995_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10784_ _06087_ VGND VGND VPWR VPWR _02110_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15311_ _02809_ VGND VGND VPWR VPWR _02810_ sky130_fd_sc_hd__clkbuf_8
X_12523_ net1965 _05735_ _07048_ VGND VGND VPWR VPWR _07083_ sky130_fd_sc_hd__mux2_1
X_16291_ CPU.registerFile\[14\]\[26\] CPU.registerFile\[10\]\[26\] _02849_ VGND VGND
+ VPWR VPWR _03764_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18030_ net1203 _02310_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_12454_ _07046_ VGND VGND VPWR VPWR _01361_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11405_ _06417_ VGND VGND VPWR VPWR _01819_ sky130_fd_sc_hd__clkbuf_1
X_12385_ _05426_ net2153 _06976_ VGND VGND VPWR VPWR _07010_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14124_ _08391_ VGND VGND VPWR VPWR _01470_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11336_ _06380_ VGND VGND VPWR VPWR _01851_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14037__314 clknet_1_0__leaf__08364_ VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__inv_2
X_11267_ CPU.registerFile\[9\]\[13\] _05708_ _06335_ VGND VGND VPWR VPWR _06344_ sky130_fd_sc_hd__mux2_1
X_13006_ CPU.registerFile\[9\]\[3\] _07283_ _07445_ _07272_ _07285_ VGND VGND VPWR
+ VPWR _07446_ sky130_fd_sc_hd__o221a_1
X_10218_ net2235 _05721_ _05713_ VGND VGND VPWR VPWR _05722_ sky130_fd_sc_hd__mux2_1
X_12768__218 clknet_1_0__leaf__07224_ VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__inv_2
X_11198_ _06307_ VGND VGND VPWR VPWR _01916_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_118_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14685__790 clknet_1_0__leaf__02684_ VGND VGND VPWR VPWR net822 sky130_fd_sc_hd__inv_2
X_17814_ net1003 _02098_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_10149_ _04713_ VGND VGND VPWR VPWR _05675_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_128_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17745_ net934 _02029_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13908_ _07330_ _08320_ VGND VGND VPWR VPWR _08321_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_18_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17676_ net865 _01964_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_141_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13839_ CPU.registerFile\[23\]\[28\] _07276_ _07618_ CPU.registerFile\[19\]\[28\]
+ _07278_ VGND VGND VPWR VPWR _08254_ sky130_fd_sc_hd__o221a_1
XFILLER_0_9_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14083__356 clknet_1_1__leaf__08368_ VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__inv_2
XFILLER_0_85_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_904 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15509_ _08397_ _02998_ _03003_ _08407_ VGND VGND VPWR VPWR _03004_ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16489_ CPU.registerFile\[26\]\[31\] _02861_ VGND VGND VPWR VPWR _03957_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09030_ CPU.cycles\[27\] _04687_ _04743_ _04708_ _04745_ VGND VGND VPWR VPWR _04746_
+ sky130_fd_sc_hd__a221o_1
X_18228_ net69 _02508_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_795 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18159_ clknet_leaf_29_clk _02439_ VGND VGND VPWR VPWR CPU.aluIn1\[25\] sky130_fd_sc_hd__dfxtp_2
Xhold302 _01493_ VGND VGND VPWR VPWR net1543 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold313 CPU.registerFile\[5\]\[6\] VGND VGND VPWR VPWR net1554 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold324 per_uart.uart0.rxd_reg\[4\] VGND VGND VPWR VPWR net1565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 CPU.registerFile\[5\]\[15\] VGND VGND VPWR VPWR net1576 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold346 per_uart.uart0.txd_reg\[6\] VGND VGND VPWR VPWR net1587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 CPU.registerFile\[2\]\[31\] VGND VGND VPWR VPWR net1598 sky130_fd_sc_hd__dlygate4sd3_1
X_14768__865 clknet_1_1__leaf__02692_ VGND VGND VPWR VPWR net897 sky130_fd_sc_hd__inv_2
X_09932_ _05556_ VGND VGND VPWR VPWR _02478_ sky130_fd_sc_hd__clkbuf_1
Xhold368 CPU.registerFile\[30\]\[24\] VGND VGND VPWR VPWR net1609 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold379 CPU.registerFile\[14\]\[31\] VGND VGND VPWR VPWR net1620 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16528__195 clknet_1_1__leaf__03964_ VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__inv_2
X_09863_ _05509_ net2046 _05491_ VGND VGND VPWR VPWR _05510_ sky130_fd_sc_hd__mux2_1
Xhold1002 CPU.registerFile\[13\]\[14\] VGND VGND VPWR VPWR net2243 sky130_fd_sc_hd__dlygate4sd3_1
X_08814_ _04528_ _04532_ _04533_ _04530_ VGND VGND VPWR VPWR _04534_ sky130_fd_sc_hd__o211ai_2
Xhold1013 CPU.registerFile\[31\]\[24\] VGND VGND VPWR VPWR net2254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1024 CPU.registerFile\[27\]\[12\] VGND VGND VPWR VPWR net2265 sky130_fd_sc_hd__dlygate4sd3_1
X_09794_ net2034 _05066_ _05463_ VGND VGND VPWR VPWR _05468_ sky130_fd_sc_hd__mux2_1
Xhold1035 CPU.registerFile\[25\]\[23\] VGND VGND VPWR VPWR net2276 sky130_fd_sc_hd__dlygate4sd3_1
X_16647__91 clknet_1_0__leaf__03989_ VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__inv_2
Xhold1046 CPU.registerFile\[21\]\[3\] VGND VGND VPWR VPWR net2287 sky130_fd_sc_hd__dlygate4sd3_1
X_08745_ _04464_ _04235_ VGND VGND VPWR VPWR _04465_ sky130_fd_sc_hd__or2_1
Xhold1057 CPU.registerFile\[6\]\[10\] VGND VGND VPWR VPWR net2298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1068 CPU.registerFile\[22\]\[28\] VGND VGND VPWR VPWR net2309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1079 CPU.registerFile\[9\]\[22\] VGND VGND VPWR VPWR net2320 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_208 _07914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08676_ _04395_ _04259_ VGND VGND VPWR VPWR _04396_ sky130_fd_sc_hd__nor2_1
XANTENNA_219 clknet_2_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_643 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09228_ _04938_ VGND VGND VPWR VPWR _04939_ sky130_fd_sc_hd__buf_4
XFILLER_0_122_907 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09159_ CPU.PC\[2\] _04870_ VGND VGND VPWR VPWR _04871_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12170_ _06861_ VGND VGND VPWR VPWR _06862_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11121_ net2156 _05698_ _06263_ VGND VGND VPWR VPWR _06267_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold880 CPU.registerFile\[20\]\[24\] VGND VGND VPWR VPWR net2121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 CPU.registerFile\[26\]\[30\] VGND VGND VPWR VPWR net2132 sky130_fd_sc_hd__dlygate4sd3_1
X_11052_ net2031 _05698_ _06226_ VGND VGND VPWR VPWR _06230_ sky130_fd_sc_hd__mux2_1
X_10003_ _04666_ _05594_ VGND VGND VPWR VPWR _05595_ sky130_fd_sc_hd__nor2_2
X_15860_ CPU.registerFile\[27\]\[13\] CPU.registerFile\[31\]\[13\] _03050_ VGND VGND
+ VPWR VPWR _03346_ sky130_fd_sc_hd__mux2_1
X_15791_ CPU.registerFile\[29\]\[11\] _02800_ VGND VGND VPWR VPWR _03279_ sky130_fd_sc_hd__or2_1
X_17530_ net719 _01818_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_11954_ CPU.registerFile\[11\]\[1\] _05733_ _06710_ VGND VGND VPWR VPWR _06744_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15234__143 clknet_1_1__leaf__02754_ VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__inv_2
X_10905_ net1715 _05687_ _06143_ VGND VGND VPWR VPWR _06152_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_123_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17461_ net650 _01749_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[16\] sky130_fd_sc_hd__dfxtp_1
X_14673_ clknet_1_1__leaf__02675_ VGND VGND VPWR VPWR _02683_ sky130_fd_sc_hd__buf_1
X_11885_ _06707_ VGND VGND VPWR VPWR _01626_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13624_ _07638_ _08043_ _08044_ _08045_ _07554_ VGND VGND VPWR VPWR _08046_ sky130_fd_sc_hd__a221o_1
X_16412_ CPU.registerFile\[15\]\[29\] CPU.registerFile\[11\]\[29\] _02849_ VGND VGND
+ VPWR VPWR _03882_ sky130_fd_sc_hd__mux2_1
X_10836_ net1951 _05687_ _06106_ VGND VGND VPWR VPWR _06115_ sky130_fd_sc_hd__mux2_1
X_17392_ net581 _01680_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13555_ _07398_ _07977_ _07978_ VGND VGND VPWR VPWR _07979_ sky130_fd_sc_hd__o21a_1
X_16343_ CPU.registerFile\[19\]\[27\] CPU.registerFile\[23\]\[27\] _02851_ VGND VGND
+ VPWR VPWR _03815_ sky130_fd_sc_hd__mux2_1
X_10767_ _06078_ VGND VGND VPWR VPWR _02118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12506_ _07074_ VGND VGND VPWR VPWR _01337_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16274_ CPU.registerFile\[17\]\[25\] _05441_ VGND VGND VPWR VPWR _03748_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13486_ CPU.registerFile\[16\]\[17\] CPU.registerFile\[20\]\[17\] _07314_ VGND VGND
+ VPWR VPWR _07912_ sky130_fd_sc_hd__mux2_1
X_10698_ _05505_ net2134 _06034_ VGND VGND VPWR VPWR _06042_ sky130_fd_sc_hd__mux2_1
X_18013_ net1186 _02293_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_12437_ _05230_ net1879 _07035_ VGND VGND VPWR VPWR _07038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12368_ _07001_ VGND VGND VPWR VPWR _01402_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14107_ net1274 _05310_ _00000_ VGND VGND VPWR VPWR _08382_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11319_ _05511_ net1969 _06371_ VGND VGND VPWR VPWR _06372_ sky130_fd_sc_hd__mux2_1
X_15087_ _07182_ net1340 VGND VGND VPWR VPWR _02273_ sky130_fd_sc_hd__nand2_1
X_12299_ CPU.aluReg\[5\] _06959_ _06861_ VGND VGND VPWR VPWR _06960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15989_ CPU.registerFile\[22\]\[17\] _08399_ VGND VGND VPWR VPWR _03471_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08530_ CPU.aluIn1\[18\] _04249_ VGND VGND VPWR VPWR _04250_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17728_ net917 _02012_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_46_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17659_ net848 _01947_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_13948__234 clknet_1_1__leaf__07226_ VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__inv_2
XFILLER_0_148_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14976__1052 clknet_1_0__leaf__02713_ VGND VGND VPWR VPWR net1084 sky130_fd_sc_hd__inv_2
X_09013_ _04716_ _04717_ _04720_ _04729_ VGND VGND VPWR VPWR _04730_ sky130_fd_sc_hd__a211o_2
XTAP_TAPCELL_ROW_154_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_154_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_586 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold110 per_uart.uart0.enable16_counter\[12\] VGND VGND VPWR VPWR net1351 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold121 mapped_spi_ram.cmd_addr\[3\] VGND VGND VPWR VPWR net1362 sky130_fd_sc_hd__dlygate4sd3_1
X_14356__494 clknet_1_0__leaf__08468_ VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__inv_2
Xhold132 mapped_spi_ram.cmd_addr\[2\] VGND VGND VPWR VPWR net1373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 mapped_spi_flash.cmd_addr\[6\] VGND VGND VPWR VPWR net1384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 mapped_spi_flash.rcv_data\[5\] VGND VGND VPWR VPWR net1395 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 mapped_spi_ram.cmd_addr\[12\] VGND VGND VPWR VPWR net1406 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold176 _07157_ VGND VGND VPWR VPWR net1417 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold187 CPU.cycles\[26\] VGND VGND VPWR VPWR net1428 sky130_fd_sc_hd__dlygate4sd3_1
X_13994__276 clknet_1_0__leaf__08359_ VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__inv_2
Xhold198 CPU.cycles\[9\] VGND VGND VPWR VPWR net1439 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09915_ _05332_ VGND VGND VPWR VPWR _05545_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09846_ _05498_ VGND VGND VPWR VPWR _02506_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_13_Left_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ net1857 _04780_ _05452_ VGND VGND VPWR VPWR _05459_ sky130_fd_sc_hd__mux2_1
X_08728_ _04447_ _04340_ VGND VGND VPWR VPWR _04448_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_1_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08659_ CPU.aluIn1\[28\] VGND VGND VPWR VPWR _04379_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14066__340 clknet_1_1__leaf__08367_ VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__inv_2
X_14521__642 clknet_1_1__leaf__02668_ VGND VGND VPWR VPWR net674 sky130_fd_sc_hd__inv_2
X_11670_ mapped_spi_ram.rcv_data\[23\] _06575_ _06586_ _06581_ VGND VGND VPWR VPWR
+ _01719_ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10621_ _05969_ VGND VGND VPWR VPWR _05994_ sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_22_Left_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13340_ _07260_ _07769_ VGND VGND VPWR VPWR _07770_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10552_ _05823_ _05949_ VGND VGND VPWR VPWR _05950_ sky130_fd_sc_hd__nand2_2
XFILLER_0_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14439__569 clknet_1_0__leaf__02659_ VGND VGND VPWR VPWR net601 sky130_fd_sc_hd__inv_2
XFILLER_0_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13271_ _07397_ _07695_ _07702_ _07703_ VGND VGND VPWR VPWR _07704_ sky130_fd_sc_hd__a31o_1
XFILLER_0_106_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10483_ _04510_ _04549_ VGND VGND VPWR VPWR _05893_ sky130_fd_sc_hd__nand2_1
X_12222_ CPU.aluIn1\[23\] _06900_ _06894_ VGND VGND VPWR VPWR _06901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12153_ _06849_ VGND VGND VPWR VPWR _01499_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11104_ net1571 _05681_ _06252_ VGND VGND VPWR VPWR _06258_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16961_ net256 _01287_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_12084_ _05359_ net1988 _06805_ VGND VGND VPWR VPWR _06813_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_31_Left_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11035_ net2140 _05681_ _06215_ VGND VGND VPWR VPWR _06221_ sky130_fd_sc_hd__mux2_1
X_15912_ _02936_ _03389_ _03396_ _02934_ VGND VGND VPWR VPWR _03397_ sky130_fd_sc_hd__o211a_1
X_16892_ per_uart.uart0.rx_bitcount\[2\] per_uart.uart0.rx_bitcount\[1\] per_uart.uart0.rx_bitcount\[0\]
+ _04137_ per_uart.uart0.rx_bitcount\[3\] VGND VGND VPWR VPWR _04172_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_125_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14905__989 clknet_1_1__leaf__02705_ VGND VGND VPWR VPWR net1021 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_125_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15843_ _02948_ _03326_ _03329_ VGND VGND VPWR VPWR _03330_ sky130_fd_sc_hd__or3_2
X_16626__72 clknet_1_0__leaf__03971_ VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__inv_2
X_14604__717 clknet_1_0__leaf__02676_ VGND VGND VPWR VPWR net749 sky130_fd_sc_hd__inv_2
XFILLER_0_59_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15774_ _03258_ _03262_ _02810_ VGND VGND VPWR VPWR _03263_ sky130_fd_sc_hd__a21o_1
X_12986_ CPU.registerFile\[18\]\[3\] CPU.registerFile\[22\]\[3\] _07240_ VGND VGND
+ VPWR VPWR _07426_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17513_ net702 _01801_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_11937_ _06735_ VGND VGND VPWR VPWR _01602_ sky130_fd_sc_hd__clkbuf_1
X_14797__891 clknet_1_0__leaf__02695_ VGND VGND VPWR VPWR net923 sky130_fd_sc_hd__inv_2
X_16641__86 clknet_1_0__leaf__03988_ VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__inv_2
X_17444_ net633 _01732_ VGND VGND VPWR VPWR mapped_spi_ram.snd_bitcount\[5\] sky130_fd_sc_hd__dfxtp_1
X_11868_ CPU.registerFile\[10\]\[10\] _05715_ _06697_ VGND VGND VPWR VPWR _06699_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10819_ _06105_ VGND VGND VPWR VPWR _06106_ sky130_fd_sc_hd__buf_4
X_13607_ CPU.registerFile\[30\]\[21\] CPU.registerFile\[26\]\[21\] _04936_ VGND VGND
+ VPWR VPWR _08029_ sky130_fd_sc_hd__mux2_1
X_17375_ net564 _01663_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11799_ _06662_ VGND VGND VPWR VPWR _01667_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_41_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16326_ CPU.registerFile\[14\]\[27\] _02826_ _02770_ VGND VGND VPWR VPWR _03798_
+ sky130_fd_sc_hd__o21a_1
X_13538_ CPU.registerFile\[5\]\[19\] CPU.registerFile\[4\]\[19\] _07577_ VGND VGND
+ VPWR VPWR _07962_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16257_ CPU.registerFile\[14\]\[25\] CPU.registerFile\[10\]\[25\] _02761_ VGND VGND
+ VPWR VPWR _03731_ sky130_fd_sc_hd__mux2_1
X_13469_ CPU.registerFile\[29\]\[17\] _07382_ _07383_ CPU.registerFile\[25\]\[17\]
+ _07570_ VGND VGND VPWR VPWR _07895_ sky130_fd_sc_hd__o221a_1
XFILLER_0_153_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650__759 clknet_1_1__leaf__02680_ VGND VGND VPWR VPWR net791 sky130_fd_sc_hd__inv_2
XFILLER_0_71_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15208_ clknet_1_1__leaf__02749_ VGND VGND VPWR VPWR _02752_ sky130_fd_sc_hd__buf_1
X_16188_ _02935_ _03657_ _03664_ _02993_ VGND VGND VPWR VPWR _03665_ sky130_fd_sc_hd__a31o_1
XFILLER_0_112_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09700_ CPU.aluIn1\[2\] net1292 VGND VGND VPWR VPWR _05391_ sky130_fd_sc_hd__or2_1
XFILLER_0_156_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09631_ _05321_ _05322_ _05323_ _05324_ _04773_ VGND VGND VPWR VPWR _05325_ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_52_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09562_ CPU.PC\[6\] _04918_ CPU.PC\[7\] VGND VGND VPWR VPWR _05258_ sky130_fd_sc_hd__a21oi_1
X_08513_ CPU.rs2\[25\] _04201_ _04206_ VGND VGND VPWR VPWR _04233_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09493_ _04758_ _05191_ _05112_ VGND VGND VPWR VPWR _05192_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_156_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09829_ net2191 _05448_ _05451_ VGND VGND VPWR VPWR _05486_ sky130_fd_sc_hd__mux2_1
X_12840_ _07238_ VGND VGND VPWR VPWR _07283_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_87_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ mapped_spi_ram.rcv_data\[0\] _06574_ _06615_ _06607_ VGND VGND VPWR VPWR
+ _01696_ sky130_fd_sc_hd__o211a_1
X_15490_ CPU.registerFile\[20\]\[3\] CPU.registerFile\[21\]\[3\] _08395_ VGND VGND
+ VPWR VPWR _02986_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11653_ _06576_ VGND VGND VPWR VPWR _06577_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_153_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10604_ net1324 _05981_ VGND VGND VPWR VPWR _05985_ sky130_fd_sc_hd__or2_1
X_17160_ net384 _01448_ VGND VGND VPWR VPWR CPU.aluReg\[24\] sky130_fd_sc_hd__dfxtp_1
X_11584_ net1406 _06517_ _06509_ _06527_ VGND VGND VPWR VPWR _06528_ sky130_fd_sc_hd__a211o_1
XFILLER_0_153_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13323_ CPU.registerFile\[15\]\[12\] _07276_ _07277_ CPU.registerFile\[11\]\[12\]
+ _07278_ VGND VGND VPWR VPWR _07754_ sky130_fd_sc_hd__o221a_1
X_16111_ CPU.registerFile\[31\]\[20\] _03072_ VGND VGND VPWR VPWR _03590_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10535_ net1367 _05892_ _05935_ _05936_ VGND VGND VPWR VPWR _02207_ sky130_fd_sc_hd__o211a_1
X_17091_ net349 _01413_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_14372__509 clknet_1_1__leaf__02652_ VGND VGND VPWR VPWR net541 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_118_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_118_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16042_ CPU.registerFile\[16\]\[18\] _02831_ _02834_ CPU.registerFile\[17\]\[18\]
+ _02854_ VGND VGND VPWR VPWR _03523_ sky130_fd_sc_hd__o221a_1
X_13254_ _07683_ _07686_ _07584_ VGND VGND VPWR VPWR _07687_ sky130_fd_sc_hd__a21oi_4
X_10466_ net1377 _05850_ _05851_ _05878_ VGND VGND VPWR VPWR _05879_ sky130_fd_sc_hd__a211o_1
Xclkbuf_1_1__f__02680_ clknet_0__02680_ VGND VGND VPWR VPWR clknet_1_1__leaf__02680_
+ sky130_fd_sc_hd__clkbuf_16
X_12205_ net2527 _06887_ _06862_ VGND VGND VPWR VPWR _06888_ sky130_fd_sc_hd__mux2_1
X_13185_ CPU.registerFile\[14\]\[8\] CPU.registerFile\[10\]\[8\] _04937_ VGND VGND
+ VPWR VPWR _07620_ sky130_fd_sc_hd__mux2_1
X_13977__260 clknet_1_1__leaf__08358_ VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__inv_2
X_10397_ _05826_ VGND VGND VPWR VPWR _05827_ sky130_fd_sc_hd__buf_2
X_12136_ _06840_ VGND VGND VPWR VPWR _01507_ sky130_fd_sc_hd__clkbuf_1
X_17993_ clknet_leaf_10_clk _02277_ VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_16944_ net239 _01270_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_12067_ _05170_ net1948 _06794_ VGND VGND VPWR VPWR _06804_ sky130_fd_sc_hd__mux2_1
X_11018_ _06211_ VGND VGND VPWR VPWR _02000_ sky130_fd_sc_hd__clkbuf_1
X_16875_ per_uart.uart0.rx_count16\[2\] _04156_ VGND VGND VPWR VPWR _04160_ sky130_fd_sc_hd__xnor2_1
X_14975__1051 clknet_1_0__leaf__02713_ VGND VGND VPWR VPWR net1083 sky130_fd_sc_hd__inv_2
X_15826_ CPU.registerFile\[29\]\[12\] _02800_ VGND VGND VPWR VPWR _03313_ sky130_fd_sc_hd__or2_1
X_15757_ _03195_ _03242_ _03243_ _03244_ _03245_ VGND VGND VPWR VPWR _03246_ sky130_fd_sc_hd__a221o_1
XFILLER_0_158_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12969_ _07401_ _07406_ _07407_ _07409_ _07360_ VGND VGND VPWR VPWR _07410_ sky130_fd_sc_hd__a221o_1
XFILLER_0_143_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15688_ CPU.registerFile\[6\]\[8\] CPU.registerFile\[7\]\[8\] _02819_ VGND VGND VPWR
+ VPWR _03179_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_380 _07570_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_391 _07305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17427_ net616 _01715_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17358_ net547 _01646_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16309_ CPU.registerFile\[27\]\[26\] CPU.registerFile\[31\]\[26\] _02852_ VGND VGND
+ VPWR VPWR _03782_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17289_ net478 _01577_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_151_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload30 clknet_1_1__leaf__03963_ VGND VGND VPWR VPWR clkload30/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_70_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload41 clknet_1_0__leaf__02744_ VGND VGND VPWR VPWR clkload41/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload52 clknet_1_1__leaf__02709_ VGND VGND VPWR VPWR clkload52/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_141_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload63 clknet_1_1__leaf__02691_ VGND VGND VPWR VPWR clkload63/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_24_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload74 clknet_1_0__leaf__02672_ VGND VGND VPWR VPWR clkload74/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload85 clknet_1_1__leaf__02659_ VGND VGND VPWR VPWR clkload85/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload96 clknet_1_0__leaf__08462_ VGND VGND VPWR VPWR clkload96/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_54_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08993_ _04216_ _04710_ _04655_ VGND VGND VPWR VPWR _04711_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_149_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14468__595 clknet_1_0__leaf__02662_ VGND VGND VPWR VPWR net627 sky130_fd_sc_hd__inv_2
XFILLER_0_97_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09614_ mapped_spi_ram.rcv_data\[13\] _04688_ _04709_ mapped_spi_flash.rcv_data\[13\]
+ VGND VGND VPWR VPWR _05308_ sky130_fd_sc_hd__a22o_4
X_09545_ _04315_ _04683_ VGND VGND VPWR VPWR _05242_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_69_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09476_ CPU.PC\[11\] _04921_ VGND VGND VPWR VPWR _05176_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload2 clknet_2_3__leaf_clk VGND VGND VPWR VPWR clkload2/Y sky130_fd_sc_hd__inv_6
XFILLER_0_33_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14633__743 clknet_1_0__leaf__02679_ VGND VGND VPWR VPWR net775 sky130_fd_sc_hd__inv_2
XFILLER_0_150_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10320_ _05497_ net2344 _05777_ VGND VGND VPWR VPWR _05781_ sky130_fd_sc_hd__mux2_1
X_17479__25 VGND VGND VPWR VPWR _17479__25/HI net25 sky130_fd_sc_hd__conb_1
X_10251_ _05497_ net2118 _05740_ VGND VGND VPWR VPWR _05744_ sky130_fd_sc_hd__mux2_1
X_10182_ _05697_ VGND VGND VPWR VPWR _02337_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13941_ _07334_ _08342_ _08345_ _08352_ _07766_ VGND VGND VPWR VPWR _08353_ sky130_fd_sc_hd__o311a_1
X_16660_ _03990_ VGND VGND VPWR VPWR _03991_ sky130_fd_sc_hd__buf_2
X_13872_ CPU.registerFile\[13\]\[29\] _07282_ _08285_ VGND VGND VPWR VPWR _08286_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_69_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15611_ CPU.registerFile\[2\]\[6\] _02821_ _02822_ CPU.registerFile\[3\]\[6\] _05070_
+ VGND VGND VPWR VPWR _03104_ sky130_fd_sc_hd__a221o_1
X_12823_ CPU.registerFile\[7\]\[0\] _07262_ _07264_ _07265_ VGND VGND VPWR VPWR _07266_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18330_ clknet_leaf_6_clk _02610_ VGND VGND VPWR VPWR per_uart.uart0.tx_count16\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_15542_ CPU.aluIn1\[4\] _02958_ _03011_ _03036_ _02995_ VGND VGND VPWR VPWR _02418_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_96_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_141_Right_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11705_ _06515_ VGND VGND VPWR VPWR _06607_ sky130_fd_sc_hd__buf_2
X_18261_ net102 _02541_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_12685_ _07170_ _07171_ VGND VGND VPWR VPWR _00034_ sky130_fd_sc_hd__nor2_1
X_15473_ CPU.registerFile\[28\]\[3\] _05049_ VGND VGND VPWR VPWR _02969_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14716__818 clknet_1_1__leaf__02687_ VGND VGND VPWR VPWR net850 sky130_fd_sc_hd__inv_2
X_17212_ net402 _01500_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11636_ net1334 _06555_ _06563_ _06474_ VGND VGND VPWR VPWR _01730_ sky130_fd_sc_hd__o22a_1
X_18192_ net223 _02472_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_115_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17143_ net367 _01431_ VGND VGND VPWR VPWR CPU.aluReg\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11567_ _06515_ VGND VGND VPWR VPWR _06516_ sky130_fd_sc_hd__buf_2
XFILLER_0_21_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_133_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13306_ CPU.rs2\[11\] _07705_ _07721_ _07736_ _07737_ VGND VGND VPWR VPWR _01306_
+ sky130_fd_sc_hd__o221a_1
X_10518_ CPU.PC\[6\] _05867_ _05922_ _05915_ VGND VGND VPWR VPWR _05923_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_133_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold709 CPU.registerFile\[10\]\[7\] VGND VGND VPWR VPWR net1950 sky130_fd_sc_hd__dlygate4sd3_1
X_17074_ net332 _01396_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11498_ _06466_ VGND VGND VPWR VPWR _01775_ sky130_fd_sc_hd__clkbuf_1
X_16025_ _03501_ _03505_ _08410_ VGND VGND VPWR VPWR _03506_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13237_ _07475_ _07669_ _07670_ VGND VGND VPWR VPWR _07671_ sky130_fd_sc_hd__o21a_1
X_10449_ net1360 _05849_ _05864_ _05855_ VGND VGND VPWR VPWR _02221_ sky130_fd_sc_hd__o211a_1
Xclkbuf_1_1__f__02663_ clknet_0__02663_ VGND VGND VPWR VPWR clknet_1_1__leaf__02663_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_122_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__02694_ _02694_ VGND VGND VPWR VPWR clknet_0__02694_ sky130_fd_sc_hd__clkbuf_16
X_13168_ _07364_ _07602_ VGND VGND VPWR VPWR _07603_ sky130_fd_sc_hd__or2_1
Xclkbuf_0__07221_ _07221_ VGND VGND VPWR VPWR clknet_0__07221_ sky130_fd_sc_hd__clkbuf_16
X_12119_ _05008_ net2076 _06830_ VGND VGND VPWR VPWR _06832_ sky130_fd_sc_hd__mux2_1
X_17976_ net1164 _02260_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_13099_ CPU.registerFile\[16\]\[6\] CPU.registerFile\[20\]\[6\] _07240_ VGND VGND
+ VPWR VPWR _07536_ sky130_fd_sc_hd__mux2_1
X_16858_ _04147_ VGND VGND VPWR VPWR _02623_ sky130_fd_sc_hd__clkbuf_1
X_15809_ _02936_ _03289_ _03296_ _02934_ VGND VGND VPWR VPWR _03297_ sky130_fd_sc_hd__o211a_1
X_16789_ _04096_ _04100_ _05815_ VGND VGND VPWR VPWR _02601_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_153_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09330_ _04445_ _05036_ VGND VGND VPWR VPWR _05037_ sky130_fd_sc_hd__xor2_1
XFILLER_0_48_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09261_ _04970_ VGND VGND VPWR VPWR _04971_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_157_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_579 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09192_ _04837_ _04902_ _04903_ VGND VGND VPWR VPWR _04904_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__08468_ _08468_ VGND VGND VPWR VPWR clknet_0__08468_ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f__08368_ clknet_0__08368_ VGND VGND VPWR VPWR clknet_1_1__leaf__08368_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08976_ _04492_ _04686_ _04694_ VGND VGND VPWR VPWR _04695_ sky130_fd_sc_hd__a21o_1
X_14214__390 clknet_1_1__leaf__08431_ VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__inv_2
Xhold69 _06620_ VGND VGND VPWR VPWR net1310 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__02752_ clknet_0__02752_ VGND VGND VPWR VPWR clknet_1_0__leaf__02752_
+ sky130_fd_sc_hd__clkbuf_16
X_15037__1108 clknet_1_0__leaf__02718_ VGND VGND VPWR VPWR net1140 sky130_fd_sc_hd__inv_2
X_16497__167 clknet_1_0__leaf__02756_ VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_84_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_84_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__02683_ clknet_0__02683_ VGND VGND VPWR VPWR clknet_1_0__leaf__02683_
+ sky130_fd_sc_hd__clkbuf_16
X_09528_ CPU.PC\[9\] _04920_ VGND VGND VPWR VPWR _05226_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09459_ _04431_ _05159_ _04400_ _04433_ VGND VGND VPWR VPWR _05160_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_47_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12470_ _07055_ VGND VGND VPWR VPWR _01354_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11421_ _05545_ net2177 _06419_ VGND VGND VPWR VPWR _06426_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14140_ _05405_ VGND VGND VPWR VPWR _08403_ sky130_fd_sc_hd__buf_4
X_11352_ _05545_ net2493 _06382_ VGND VGND VPWR VPWR _06389_ sky130_fd_sc_hd__mux2_1
X_14974__1050 clknet_1_0__leaf__02713_ VGND VGND VPWR VPWR net1082 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_115_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10303_ _05549_ net2245 _05762_ VGND VGND VPWR VPWR _05771_ sky130_fd_sc_hd__mux2_1
X_11283_ _06352_ VGND VGND VPWR VPWR _01876_ sky130_fd_sc_hd__clkbuf_1
X_13022_ CPU.registerFile\[6\]\[4\] CPU.registerFile\[7\]\[4\] _07371_ VGND VGND VPWR
+ VPWR _07461_ sky130_fd_sc_hd__mux2_1
X_10234_ _05732_ VGND VGND VPWR VPWR _02320_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_5_Left_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17830_ net1019 _02114_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_10165_ net1821 _05685_ _05671_ VGND VGND VPWR VPWR _05686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17761_ net950 _02045_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_14973_ clknet_1_1__leaf__02708_ VGND VGND VPWR VPWR _02713_ sky130_fd_sc_hd__buf_1
X_10096_ _05645_ VGND VGND VPWR VPWR _02371_ sky130_fd_sc_hd__clkbuf_1
X_16712_ _04001_ _05218_ VGND VGND VPWR VPWR _04036_ sky130_fd_sc_hd__nand2_1
X_13924_ CPU.registerFile\[21\]\[31\] _07347_ _07429_ CPU.registerFile\[17\]\[31\]
+ _07349_ VGND VGND VPWR VPWR _08336_ sky130_fd_sc_hd__o221a_1
X_17692_ net881 _01980_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13855_ _07801_ _08266_ _08267_ _08268_ _07555_ VGND VGND VPWR VPWR _08269_ sky130_fd_sc_hd__a221o_1
XFILLER_0_69_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12806_ _04970_ VGND VGND VPWR VPWR _07249_ sky130_fd_sc_hd__buf_4
X_10998_ _06178_ VGND VGND VPWR VPWR _06201_ sky130_fd_sc_hd__clkbuf_4
X_13786_ _07231_ _08199_ _08202_ VGND VGND VPWR VPWR _08203_ sky130_fd_sc_hd__or3_1
XFILLER_0_69_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18313_ clknet_leaf_16_clk _02593_ VGND VGND VPWR VPWR CPU.PC\[13\] sky130_fd_sc_hd__dfxtp_1
X_15525_ _03015_ _03016_ _03018_ _03019_ VGND VGND VPWR VPWR _03020_ sky130_fd_sc_hd__o211a_1
X_14304__447 clknet_1_1__leaf__08463_ VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__inv_2
X_12737_ _07214_ VGND VGND VPWR VPWR _01260_ sky130_fd_sc_hd__clkbuf_1
X_16929__9 clknet_1_1__leaf__07220_ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__inv_2
XFILLER_0_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18244_ net85 _02524_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_15456_ CPU.registerFile\[22\]\[2\] CPU.registerFile\[23\]\[2\] _02829_ VGND VGND
+ VPWR VPWR _02953_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12668_ _07160_ net1380 VGND VGND VPWR VPWR _00027_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14407_ clknet_1_0__leaf__02653_ VGND VGND VPWR VPWR _02657_ sky130_fd_sc_hd__buf_1
X_18175_ net206 _02455_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_11619_ mapped_spi_ram.snd_bitcount\[2\] mapped_spi_ram.snd_bitcount\[1\] mapped_spi_ram.snd_bitcount\[0\]
+ VGND VGND VPWR VPWR _06549_ sky130_fd_sc_hd__or3_1
X_15387_ _02796_ VGND VGND VPWR VPWR _02885_ sky130_fd_sc_hd__buf_4
XFILLER_0_41_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12599_ net1329 _05822_ _05942_ VGND VGND VPWR VPWR _00006_ sky130_fd_sc_hd__o21a_1
XFILLER_0_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17126_ clknet_leaf_20_clk _00029_ VGND VGND VPWR VPWR CPU.cycles\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold506 per_uart.d_in_uart\[7\] VGND VGND VPWR VPWR net1747 sky130_fd_sc_hd__dlygate4sd3_1
Xhold517 CPU.registerFile\[22\]\[21\] VGND VGND VPWR VPWR net1758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold528 CPU.registerFile\[13\]\[31\] VGND VGND VPWR VPWR net1769 sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 CPU.registerFile\[3\]\[1\] VGND VGND VPWR VPWR net1780 sky130_fd_sc_hd__dlygate4sd3_1
X_17057_ net315 _01379_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[19\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__02715_ clknet_0__02715_ VGND VGND VPWR VPWR clknet_1_1__leaf__02715_
+ sky130_fd_sc_hd__clkbuf_16
X_14269_ _04485_ _06872_ _08447_ VGND VGND VPWR VPWR _08448_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16008_ CPU.registerFile\[27\]\[17\] _02928_ _02910_ VGND VGND VPWR VPWR _03490_
+ sky130_fd_sc_hd__o21a_1
Xclkbuf_0__02746_ _02746_ VGND VGND VPWR VPWR clknet_0__02746_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_21_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08830_ _04548_ _04510_ _04549_ VGND VGND VPWR VPWR _04550_ sky130_fd_sc_hd__a21bo_1
Xclkbuf_0__02677_ _02677_ VGND VGND VPWR VPWR clknet_0__02677_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_148_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14350__489 clknet_1_1__leaf__08467_ VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__inv_2
Xhold1206 CPU.registerFile\[11\]\[8\] VGND VGND VPWR VPWR net2447 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1217 CPU.registerFile\[8\]\[12\] VGND VGND VPWR VPWR net2458 sky130_fd_sc_hd__dlygate4sd3_1
X_08761_ _04370_ _04478_ _04480_ VGND VGND VPWR VPWR _04481_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_146_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1228 CPU.registerFile\[16\]\[12\] VGND VGND VPWR VPWR net2469 sky130_fd_sc_hd__dlygate4sd3_1
X_17959_ net1147 _02243_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[4\] sky130_fd_sc_hd__dfxtp_1
Xhold1239 CPU.registerFile\[2\]\[12\] VGND VGND VPWR VPWR net2480 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08692_ CPU.aluIn1\[0\] VGND VGND VPWR VPWR _04412_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_49_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09313_ _05017_ _05018_ _05020_ _04773_ VGND VGND VPWR VPWR _05021_ sky130_fd_sc_hd__o31a_1
XFILLER_0_48_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09244_ _04915_ VGND VGND VPWR VPWR _04955_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_62_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14060__335 clknet_1_1__leaf__08366_ VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_32_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09175_ _04860_ _04885_ _04886_ VGND VGND VPWR VPWR _04887_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14745__844 clknet_1_1__leaf__02690_ VGND VGND VPWR VPWR net876 sky130_fd_sc_hd__inv_2
X_08959_ _04677_ VGND VGND VPWR VPWR _04678_ sky130_fd_sc_hd__clkbuf_4
X_16505__174 clknet_1_1__leaf__03962_ VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__inv_2
X_11970_ _04762_ net1764 _06747_ VGND VGND VPWR VPWR _06753_ sky130_fd_sc_hd__mux2_1
X_10921_ _06160_ VGND VGND VPWR VPWR _02046_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10852_ _06123_ VGND VGND VPWR VPWR _02078_ sky130_fd_sc_hd__clkbuf_1
X_13640_ CPU.registerFile\[23\]\[22\] _07244_ _07429_ CPU.registerFile\[19\]\[22\]
+ _07820_ VGND VGND VPWR VPWR _08061_ sky130_fd_sc_hd__o221a_1
Xclkbuf_1_0__f__02666_ clknet_0__02666_ VGND VGND VPWR VPWR clknet_1_0__leaf__02666_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_66_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_866 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10783_ _05522_ net1852 _06081_ VGND VGND VPWR VPWR _06087_ sky130_fd_sc_hd__mux2_1
X_13571_ CPU.registerFile\[19\]\[20\] _07618_ _07993_ _07417_ _07253_ VGND VGND VPWR
+ VPWR _07994_ sky130_fd_sc_hd__o221a_1
XFILLER_0_82_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15310_ _05010_ VGND VGND VPWR VPWR _02809_ sky130_fd_sc_hd__buf_6
X_12522_ _07082_ VGND VGND VPWR VPWR _01329_ sky130_fd_sc_hd__clkbuf_1
X_16290_ CPU.aluIn1\[25\] _07358_ _03763_ _03632_ VGND VGND VPWR VPWR _02439_ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14791__886 clknet_1_0__leaf__02694_ VGND VGND VPWR VPWR net918 sky130_fd_sc_hd__inv_2
XFILLER_0_152_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15241_ clknet_1_1__leaf__02749_ VGND VGND VPWR VPWR _02755_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_10_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12453_ _05426_ net2012 _07012_ VGND VGND VPWR VPWR _07046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14490__614 clknet_1_0__leaf__02665_ VGND VGND VPWR VPWR net646 sky130_fd_sc_hd__inv_2
XFILLER_0_151_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11404_ _05528_ net1949 _06408_ VGND VGND VPWR VPWR _06417_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12384_ _07009_ VGND VGND VPWR VPWR _01394_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14123_ _04208_ _05152_ _08387_ VGND VGND VPWR VPWR _08391_ sky130_fd_sc_hd__mux2_1
X_11335_ _05528_ net1883 _06371_ VGND VGND VPWR VPWR _06380_ sky130_fd_sc_hd__mux2_1
X_14828__919 clknet_1_1__leaf__02698_ VGND VGND VPWR VPWR net951 sky130_fd_sc_hd__inv_2
X_11266_ _06343_ VGND VGND VPWR VPWR _01884_ sky130_fd_sc_hd__clkbuf_1
X_14054_ clknet_1_1__leaf__08363_ VGND VGND VPWR VPWR _08366_ sky130_fd_sc_hd__buf_1
XFILLER_0_120_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10217_ _05272_ VGND VGND VPWR VPWR _05721_ sky130_fd_sc_hd__clkbuf_4
X_13005_ CPU.registerFile\[8\]\[3\] CPU.registerFile\[12\]\[3\] _07339_ VGND VGND
+ VPWR VPWR _07445_ sky130_fd_sc_hd__mux2_1
X_14230__405 clknet_1_1__leaf__08432_ VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__inv_2
XFILLER_0_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11197_ _05526_ net2090 _06299_ VGND VGND VPWR VPWR _06307_ sky130_fd_sc_hd__mux2_1
X_17813_ net1002 _02097_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_10148_ _05674_ VGND VGND VPWR VPWR _02348_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_128_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17744_ net933 _02028_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_10079_ _05636_ VGND VGND VPWR VPWR _02379_ sky130_fd_sc_hd__clkbuf_1
X_13907_ CPU.registerFile\[28\]\[30\] CPU.registerFile\[24\]\[30\] _07352_ VGND VGND
+ VPWR VPWR _08320_ sky130_fd_sc_hd__mux2_1
X_17675_ net864 _01963_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_59_Left_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_141_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_141_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13838_ CPU.registerFile\[18\]\[28\] CPU.registerFile\[22\]\[28\] _07648_ VGND VGND
+ VPWR VPWR _08253_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15211__122 clknet_1_1__leaf__02752_ VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__inv_2
X_13769_ CPU.registerFile\[21\]\[26\] _07403_ _07404_ CPU.registerFile\[17\]\[26\]
+ _07250_ VGND VGND VPWR VPWR _08186_ sky130_fd_sc_hd__o221a_1
XFILLER_0_85_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15508_ _02914_ _03000_ _03002_ _02965_ VGND VGND VPWR VPWR _03003_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_44_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16488_ CPU.registerFile\[28\]\[31\] CPU.registerFile\[24\]\[31\] _02761_ VGND VGND
+ VPWR VPWR _03956_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18227_ net68 _02507_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15439_ _05361_ VGND VGND VPWR VPWR _02936_ sky130_fd_sc_hd__buf_2
XFILLER_0_115_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18158_ clknet_leaf_29_clk _02438_ VGND VGND VPWR VPWR CPU.aluIn1\[24\] sky130_fd_sc_hd__dfxtp_2
XPHY_EDGE_ROW_68_Left_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold303 CPU.PC\[18\] VGND VGND VPWR VPWR net1544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 CPU.registerFile\[6\]\[1\] VGND VGND VPWR VPWR net1555 sky130_fd_sc_hd__dlygate4sd3_1
X_17109_ clknet_leaf_23_clk _00042_ VGND VGND VPWR VPWR CPU.cycles\[5\] sky130_fd_sc_hd__dfxtp_1
X_15036__1107 clknet_1_0__leaf__02718_ VGND VGND VPWR VPWR net1139 sky130_fd_sc_hd__inv_2
XFILLER_0_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold325 _04144_ VGND VGND VPWR VPWR net1566 sky130_fd_sc_hd__dlygate4sd3_1
X_18089_ net152 _02369_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold336 CPU.registerFile\[6\]\[31\] VGND VGND VPWR VPWR net1577 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold347 CPU.PC\[16\] VGND VGND VPWR VPWR net1588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 CPU.registerFile\[5\]\[26\] VGND VGND VPWR VPWR net1599 sky130_fd_sc_hd__dlygate4sd3_1
X_09931_ _05555_ net1716 _05490_ VGND VGND VPWR VPWR _05556_ sky130_fd_sc_hd__mux2_1
Xhold369 mapped_spi_ram.rcv_data\[19\] VGND VGND VPWR VPWR net1610 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09862_ _04957_ VGND VGND VPWR VPWR _05509_ sky130_fd_sc_hd__buf_4
XFILLER_0_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08813_ CPU.aluIn1\[3\] _04521_ VGND VGND VPWR VPWR _04533_ sky130_fd_sc_hd__nand2_1
Xhold1003 CPU.registerFile\[21\]\[18\] VGND VGND VPWR VPWR net2244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1014 CPU.registerFile\[25\]\[30\] VGND VGND VPWR VPWR net2255 sky130_fd_sc_hd__dlygate4sd3_1
X_09793_ _05467_ VGND VGND VPWR VPWR _02528_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1025 CPU.registerFile\[2\]\[10\] VGND VGND VPWR VPWR net2266 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1036 CPU.registerFile\[31\]\[27\] VGND VGND VPWR VPWR net2277 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1047 CPU.registerFile\[31\]\[15\] VGND VGND VPWR VPWR net2288 sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ CPU.aluIn1\[24\] VGND VGND VPWR VPWR _04464_ sky130_fd_sc_hd__inv_2
Xhold1058 CPU.registerFile\[16\]\[11\] VGND VGND VPWR VPWR net2299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1069 CPU.registerFile\[15\]\[26\] VGND VGND VPWR VPWR net2310 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_77_Left_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08675_ CPU.aluIn1\[13\] VGND VGND VPWR VPWR _04395_ sky130_fd_sc_hd__inv_2
XANTENNA_209 _07914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09227_ _04937_ VGND VGND VPWR VPWR _04938_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_86_Left_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09158_ CPU.instr\[3\] CPU.Iimm\[2\] _04664_ _04830_ VGND VGND VPWR VPWR _04870_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09089_ _04461_ _04457_ _04459_ VGND VGND VPWR VPWR _04801_ sky130_fd_sc_hd__nor3_1
XFILLER_0_4_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11120_ _06266_ VGND VGND VPWR VPWR _01953_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_92_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold870 CPU.registerFile\[21\]\[21\] VGND VGND VPWR VPWR net2111 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold881 CPU.registerFile\[23\]\[30\] VGND VGND VPWR VPWR net2122 sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ _06229_ VGND VGND VPWR VPWR _01985_ sky130_fd_sc_hd__clkbuf_1
Xhold892 CPU.registerFile\[30\]\[11\] VGND VGND VPWR VPWR net2133 sky130_fd_sc_hd__dlygate4sd3_1
X_14333__473 clknet_1_0__leaf__08466_ VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__inv_2
XFILLER_0_101_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10002_ _04660_ _04661_ VGND VGND VPWR VPWR _05594_ sky130_fd_sc_hd__nand2b_4
X_13971__255 clknet_1_1__leaf__08357_ VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_95_Left_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15790_ CPU.registerFile\[27\]\[11\] CPU.registerFile\[31\]\[11\] _03050_ VGND VGND
+ VPWR VPWR _03278_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11953_ _06743_ VGND VGND VPWR VPWR _01594_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10904_ _06151_ VGND VGND VPWR VPWR _02054_ sky130_fd_sc_hd__clkbuf_1
X_17460_ net649 _01748_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_123_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11884_ net2300 _05731_ _06697_ VGND VGND VPWR VPWR _06707_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__02718_ clknet_0__02718_ VGND VGND VPWR VPWR clknet_1_0__leaf__02718_
+ sky130_fd_sc_hd__clkbuf_16
X_16411_ _03195_ _03878_ _03879_ _03880_ _03245_ VGND VGND VPWR VPWR _03881_ sky130_fd_sc_hd__a221o_1
X_13623_ CPU.registerFile\[3\]\[21\] _07262_ _04938_ VGND VGND VPWR VPWR _08045_ sky130_fd_sc_hd__o21a_1
XFILLER_0_67_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10835_ _06114_ VGND VGND VPWR VPWR _02086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17391_ net580 _01679_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_24_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_109_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16342_ _05071_ _03813_ _02870_ VGND VGND VPWR VPWR _03814_ sky130_fd_sc_hd__a21o_1
X_13554_ CPU.registerFile\[29\]\[19\] _07629_ _07488_ CPU.registerFile\[25\]\[19\]
+ _04971_ VGND VGND VPWR VPWR _07978_ sky130_fd_sc_hd__o221a_1
XFILLER_0_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10766_ _05505_ net1609 _06070_ VGND VGND VPWR VPWR _06078_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12505_ net1830 _05717_ _07071_ VGND VGND VPWR VPWR _07074_ sky130_fd_sc_hd__mux2_1
X_16273_ _02810_ _03734_ _03738_ _03746_ VGND VGND VPWR VPWR _03747_ sky130_fd_sc_hd__a31o_1
X_10697_ _06041_ VGND VGND VPWR VPWR _02151_ sky130_fd_sc_hd__clkbuf_1
X_13485_ CPU.registerFile\[21\]\[17\] _07502_ _07503_ CPU.registerFile\[17\]\[17\]
+ _07300_ VGND VGND VPWR VPWR _07911_ sky130_fd_sc_hd__o221a_1
XFILLER_0_23_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18012_ net1185 _02292_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_12774__223 clknet_1_1__leaf__07225_ VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__inv_2
XFILLER_0_82_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12436_ _07037_ VGND VGND VPWR VPWR _01370_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_755 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14416__548 clknet_1_1__leaf__02657_ VGND VGND VPWR VPWR net580 sky130_fd_sc_hd__inv_2
X_12367_ _05209_ CPU.registerFile\[29\]\[10\] _06999_ VGND VGND VPWR VPWR _07001_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14106_ _08381_ VGND VGND VPWR VPWR _01462_ sky130_fd_sc_hd__clkbuf_1
X_11318_ _06359_ VGND VGND VPWR VPWR _06371_ sky130_fd_sc_hd__buf_4
X_15086_ net1339 _07181_ _02726_ VGND VGND VPWR VPWR _02730_ sky130_fd_sc_hd__a21oi_1
X_12298_ CPU.aluIn1\[5\] _06958_ _06859_ VGND VGND VPWR VPWR _06959_ sky130_fd_sc_hd__mux2_1
X_11249_ _06334_ VGND VGND VPWR VPWR _01892_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_143_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15988_ CPU.registerFile\[21\]\[17\] CPU.registerFile\[23\]\[17\] _05441_ VGND VGND
+ VPWR VPWR _03470_ sky130_fd_sc_hd__mux2_1
X_17727_ net916 _02011_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17658_ net847 _01946_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_46_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16609_ net1540 net1508 _03979_ VGND VGND VPWR VPWR _03980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17589_ net778 _01877_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[7\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_15_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_836 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14774__870 clknet_1_1__leaf__02693_ VGND VGND VPWR VPWR net902 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_158_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09012_ _04722_ _04728_ _04492_ VGND VGND VPWR VPWR _04729_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_154_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold100 per_uart.uart0.enable16_counter\[0\] VGND VGND VPWR VPWR net1341 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold111 per_uart.uart0.enable16_counter\[6\] VGND VGND VPWR VPWR net1352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 per_uart.uart0.enable16_counter\[1\] VGND VGND VPWR VPWR net1363 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold133 mapped_spi_flash.cmd_addr\[20\] VGND VGND VPWR VPWR net1374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 mapped_spi_flash.cmd_addr\[21\] VGND VGND VPWR VPWR net1385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 _02172_ VGND VGND VPWR VPWR net1396 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 mapped_spi_ram.rcv_data\[29\] VGND VGND VPWR VPWR net1407 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold177 mapped_spi_flash.state\[2\] VGND VGND VPWR VPWR net1418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 _07169_ VGND VGND VPWR VPWR net1429 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold199 per_uart.uart0.enable16_counter\[8\] VGND VGND VPWR VPWR net1440 sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ _05544_ VGND VGND VPWR VPWR _02484_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_74_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09845_ _05497_ net2068 _05491_ VGND VGND VPWR VPWR _05498_ sky130_fd_sc_hd__mux2_1
X_09776_ _05458_ VGND VGND VPWR VPWR _02536_ sky130_fd_sc_hd__clkbuf_1
X_08727_ CPU.aluIn1\[19\] _04247_ VGND VGND VPWR VPWR _04447_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ _04377_ _04223_ VGND VGND VPWR VPWR _04378_ sky130_fd_sc_hd__nor2_1
X_14857__945 clknet_1_1__leaf__02701_ VGND VGND VPWR VPWR net977 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_105_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_105_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08589_ _04308_ VGND VGND VPWR VPWR _04309_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10620_ net2467 _05983_ _05992_ _05993_ VGND VGND VPWR VPWR _02179_ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10551_ mapped_spi_flash.state\[2\] _05817_ mapped_spi_flash.state\[0\] net2 VGND
+ VGND VPWR VPWR _05949_ sky130_fd_sc_hd__o31a_1
XFILLER_0_134_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13270_ _07308_ VGND VGND VPWR VPWR _07703_ sky130_fd_sc_hd__buf_4
X_10482_ _05842_ VGND VGND VPWR VPWR _05892_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_20_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12221_ CPU.aluReg\[24\] CPU.aluReg\[22\] _06871_ VGND VGND VPWR VPWR _06900_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12152_ _05359_ net1841 _06841_ VGND VGND VPWR VPWR _06849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11103_ _06257_ VGND VGND VPWR VPWR _01961_ sky130_fd_sc_hd__clkbuf_1
X_16960_ net255 _01286_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_12083_ _06812_ VGND VGND VPWR VPWR _01532_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_9_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11034_ _06220_ VGND VGND VPWR VPWR _01993_ sky130_fd_sc_hd__clkbuf_1
X_15911_ _02948_ _03392_ _03395_ VGND VGND VPWR VPWR _03396_ sky130_fd_sc_hd__or3_2
X_16891_ net1684 VGND VGND VPWR VPWR _04171_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_125_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15842_ _02926_ _03327_ _03328_ VGND VGND VPWR VPWR _03329_ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15773_ _02914_ _03259_ _03261_ _02864_ VGND VGND VPWR VPWR _03262_ sky130_fd_sc_hd__a211o_1
X_12985_ CPU.mem_wdata\[2\] _07358_ _07396_ _07425_ _05844_ VGND VGND VPWR VPWR _01297_
+ sky130_fd_sc_hd__o221a_1
X_17512_ net701 _01800_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_736 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15035__1106 clknet_1_1__leaf__02718_ VGND VGND VPWR VPWR net1138 sky130_fd_sc_hd__inv_2
X_11936_ CPU.registerFile\[11\]\[10\] _05715_ _06733_ VGND VGND VPWR VPWR _06735_
+ sky130_fd_sc_hd__mux2_1
X_17443_ net632 _01731_ VGND VGND VPWR VPWR mapped_spi_ram.snd_bitcount\[4\] sky130_fd_sc_hd__dfxtp_1
X_11867_ _06698_ VGND VGND VPWR VPWR _01635_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13606_ CPU.registerFile\[29\]\[21\] _07772_ _07773_ CPU.registerFile\[25\]\[21\]
+ _08027_ VGND VGND VPWR VPWR _08028_ sky130_fd_sc_hd__o221a_1
X_10818_ _05631_ _05669_ VGND VGND VPWR VPWR _06105_ sky130_fd_sc_hd__nor2_4
XFILLER_0_27_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17374_ net563 _01662_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11798_ _05188_ net2308 _06661_ VGND VGND VPWR VPWR _06662_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_41_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16325_ CPU.registerFile\[10\]\[27\] _03280_ VGND VGND VPWR VPWR _03797_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13537_ _07392_ _07956_ _07960_ _07271_ VGND VGND VPWR VPWR _07961_ sky130_fd_sc_hd__o211a_2
XFILLER_0_153_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10749_ _06068_ VGND VGND VPWR VPWR _02126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16256_ CPU.aluIn1\[24\] _07358_ _03730_ _03632_ VGND VGND VPWR VPWR _02438_ sky130_fd_sc_hd__o211a_1
X_13468_ CPU.registerFile\[28\]\[17\] CPU.registerFile\[24\]\[17\] _04939_ VGND VGND
+ VPWR VPWR _07894_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_136_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12419_ _07028_ VGND VGND VPWR VPWR _01378_ sky130_fd_sc_hd__clkbuf_1
X_16187_ _05361_ _03663_ VGND VGND VPWR VPWR _03664_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13399_ CPU.registerFile\[29\]\[14\] _07556_ _07557_ CPU.registerFile\[25\]\[14\]
+ _07827_ VGND VGND VPWR VPWR _07828_ sky130_fd_sc_hd__o221a_1
XFILLER_0_10_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_4_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_155_Right_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09630_ _04311_ _04214_ _04219_ CPU.aluReg\[5\] VGND VGND VPWR VPWR _05324_ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14015__295 clknet_1_1__leaf__08361_ VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__inv_2
X_09561_ _05256_ _04883_ VGND VGND VPWR VPWR _05257_ sky130_fd_sc_hd__xor2_1
X_08512_ CPU.aluIn1\[26\] _04231_ VGND VGND VPWR VPWR _04232_ sky130_fd_sc_hd__and2_1
X_09492_ mapped_spi_ram.rcv_data\[18\] _04689_ _04691_ mapped_spi_flash.rcv_data\[18\]
+ VGND VGND VPWR VPWR _05191_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_122_Right_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09828_ _05485_ VGND VGND VPWR VPWR _02511_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_107_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09759_ _05447_ VGND VGND VPWR VPWR _05448_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_87_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14445__574 clknet_1_0__leaf__02660_ VGND VGND VPWR VPWR net606 sky130_fd_sc_hd__inv_2
X_12770_ clknet_1_1__leaf__07223_ VGND VGND VPWR VPWR _07225_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_87_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ net1473 _06576_ VGND VGND VPWR VPWR _06615_ sky130_fd_sc_hd__or2_1
X_14183__362 clknet_1_1__leaf__08428_ VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__inv_2
XFILLER_0_96_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14440_ clknet_1_1__leaf__02653_ VGND VGND VPWR VPWR _02660_ sky130_fd_sc_hd__buf_1
XFILLER_0_127_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11652_ net8 mapped_spi_ram.state\[3\] _06572_ VGND VGND VPWR VPWR _06576_ sky130_fd_sc_hd__and3_1
XFILLER_0_138_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10603_ net1324 _05983_ _05984_ _05980_ VGND VGND VPWR VPWR _02187_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11583_ _06512_ _05919_ VGND VGND VPWR VPWR _06527_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16110_ CPU.registerFile\[25\]\[20\] CPU.registerFile\[29\]\[20\] _03254_ VGND VGND
+ VPWR VPWR _03589_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13322_ CPU.registerFile\[14\]\[12\] CPU.registerFile\[10\]\[12\] _07274_ VGND VGND
+ VPWR VPWR _07753_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17090_ net348 _01412_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_10534_ _05843_ VGND VGND VPWR VPWR _05936_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16041_ CPU.registerFile\[20\]\[18\] CPU.registerFile\[21\]\[18\] _08394_ VGND VGND
+ VPWR VPWR _03522_ sky130_fd_sc_hd__mux2_1
X_10465_ _05852_ _05877_ VGND VGND VPWR VPWR _05878_ sky130_fd_sc_hd__nor2_1
X_13253_ _07653_ _07684_ _07685_ VGND VGND VPWR VPWR _07686_ sky130_fd_sc_hd__o21ai_2
X_14911__994 clknet_1_1__leaf__02706_ VGND VGND VPWR VPWR net1026 sky130_fd_sc_hd__inv_2
XFILLER_0_122_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12204_ CPU.aluIn1\[27\] _06886_ _06865_ VGND VGND VPWR VPWR _06887_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14610__722 clknet_1_0__leaf__02677_ VGND VGND VPWR VPWR net754 sky130_fd_sc_hd__inv_2
X_13184_ _07618_ VGND VGND VPWR VPWR _07619_ sky130_fd_sc_hd__buf_6
X_10396_ mapped_spi_flash.state\[2\] _05817_ _05823_ VGND VGND VPWR VPWR _05826_ sky130_fd_sc_hd__o21ai_1
X_12135_ _05170_ net2265 _06830_ VGND VGND VPWR VPWR _06840_ sky130_fd_sc_hd__mux2_1
X_17992_ clknet_leaf_10_clk net1353 VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_16943_ net238 _01269_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12066_ _06803_ VGND VGND VPWR VPWR _01540_ sky130_fd_sc_hd__clkbuf_1
X_11017_ net1626 _05731_ _06201_ VGND VGND VPWR VPWR _06211_ sky130_fd_sc_hd__mux2_1
X_14528__649 clknet_1_0__leaf__02668_ VGND VGND VPWR VPWR net681 sky130_fd_sc_hd__inv_2
X_16874_ _06030_ _04159_ VGND VGND VPWR VPWR _02627_ sky130_fd_sc_hd__nor2_1
X_15825_ CPU.registerFile\[27\]\[12\] CPU.registerFile\[31\]\[12\] _03050_ VGND VGND
+ VPWR VPWR _03312_ sky130_fd_sc_hd__mux2_1
X_15756_ _02870_ VGND VGND VPWR VPWR _03245_ sky130_fd_sc_hd__buf_4
X_12968_ _07398_ _07408_ VGND VGND VPWR VPWR _07409_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14707_ clknet_1_0__leaf__02686_ VGND VGND VPWR VPWR _02687_ sky130_fd_sc_hd__buf_1
X_11919_ CPU.registerFile\[11\]\[18\] _05698_ _06722_ VGND VGND VPWR VPWR _06726_
+ sky130_fd_sc_hd__mux2_1
X_15687_ CPU.registerFile\[1\]\[8\] _02814_ _03177_ _02816_ VGND VGND VPWR VPWR _03178_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_370 _05380_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12899_ CPU.registerFile\[9\]\[1\] _07283_ _07340_ _07272_ _07285_ VGND VGND VPWR
+ VPWR _07341_ sky130_fd_sc_hd__o221a_1
XANTENNA_381 _07621_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_392 _07318_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17426_ net615 _01714_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17357_ net546 _01645_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16308_ _03779_ _03780_ _08400_ VGND VGND VPWR VPWR _03781_ sky130_fd_sc_hd__mux2_1
X_17288_ net477 _01576_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload20 clknet_leaf_4_clk VGND VGND VPWR VPWR clkload20/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_151_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16239_ _02885_ _03711_ _03712_ _03713_ _03022_ VGND VGND VPWR VPWR _03714_ sky130_fd_sc_hd__a221o_1
Xclkload31 clknet_1_0__leaf__02755_ VGND VGND VPWR VPWR clkload31/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload42 clknet_1_1__leaf__02743_ VGND VGND VPWR VPWR clkload42/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_2_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload53 clknet_1_1__leaf__02706_ VGND VGND VPWR VPWR clkload53/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload64 clknet_1_1__leaf__02687_ VGND VGND VPWR VPWR clkload64/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_3_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload75 clknet_1_0__leaf__02671_ VGND VGND VPWR VPWR clkload75/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_2_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload86 clknet_1_1__leaf__02658_ VGND VGND VPWR VPWR clkload86/Y sky130_fd_sc_hd__clkinvlp_4
X_14886__971 clknet_1_0__leaf__02704_ VGND VGND VPWR VPWR net1003 sky130_fd_sc_hd__inv_2
Xclkload97 clknet_1_1__leaf__08435_ VGND VGND VPWR VPWR clkload97/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_54_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08992_ mapped_spi_ram.rcv_data\[5\] _04688_ _04709_ mapped_spi_flash.rcv_data\[5\]
+ VGND VGND VPWR VPWR _04710_ sky130_fd_sc_hd__a22o_2
XFILLER_0_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_149_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09613_ _05307_ VGND VGND VPWR VPWR _02556_ sky130_fd_sc_hd__clkbuf_1
X_09544_ _04920_ _05240_ VGND VGND VPWR VPWR _05241_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_69_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09475_ _04856_ _04891_ VGND VGND VPWR VPWR _05175_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload3 clknet_leaf_22_clk VGND VGND VPWR VPWR clkload3/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10250_ _05743_ VGND VGND VPWR VPWR _02315_ sky130_fd_sc_hd__clkbuf_1
X_15034__1105 clknet_1_1__leaf__02718_ VGND VGND VPWR VPWR net1137 sky130_fd_sc_hd__inv_2
XFILLER_0_30_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10181_ net2189 _05696_ _05692_ VGND VGND VPWR VPWR _05697_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13940_ _07250_ _08348_ _08349_ _08351_ _07359_ VGND VGND VPWR VPWR _08352_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_89_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15049__1116 clknet_1_0__leaf__02721_ VGND VGND VPWR VPWR net1148 sky130_fd_sc_hd__inv_2
X_13871_ CPU.registerFile\[9\]\[29\] _07618_ _08284_ _07417_ _07554_ VGND VGND VPWR
+ VPWR _08285_ sky130_fd_sc_hd__o221a_1
X_15610_ CPU.registerFile\[6\]\[6\] CPU.registerFile\[7\]\[6\] _02819_ VGND VGND VPWR
+ VPWR _03103_ sky130_fd_sc_hd__mux2_1
X_12822_ _05283_ VGND VGND VPWR VPWR _07265_ sky130_fd_sc_hd__buf_4
XFILLER_0_57_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15541_ _08411_ _03021_ _03035_ _02993_ VGND VGND VPWR VPWR _03036_ sky130_fd_sc_hd__a31o_1
XFILLER_0_97_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11704_ mapped_spi_ram.rcv_data\[9\] _06601_ VGND VGND VPWR VPWR _06606_ sky130_fd_sc_hd__or2_1
X_18260_ net101 _02540_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_15472_ CPU.registerFile\[30\]\[3\] CPU.registerFile\[26\]\[3\] _02918_ VGND VGND
+ VPWR VPWR _02968_ sky130_fd_sc_hd__mux2_1
X_12684_ net1489 _07168_ VGND VGND VPWR VPWR _07171_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17211_ net401 _01499_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_18191_ net222 _02471_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_11635_ _06499_ _06561_ _06562_ VGND VGND VPWR VPWR _06563_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17142_ net366 _01430_ VGND VGND VPWR VPWR CPU.aluReg\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11566_ _04192_ VGND VGND VPWR VPWR _06515_ sky130_fd_sc_hd__buf_4
XFILLER_0_13_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13305_ _05843_ VGND VGND VPWR VPWR _07737_ sky130_fd_sc_hd__buf_2
XFILLER_0_52_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17073_ net331 _01395_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_10517_ net1278 _04541_ _04590_ VGND VGND VPWR VPWR _05922_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_133_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14285_ clknet_1_1__leaf__08433_ VGND VGND VPWR VPWR _08462_ sky130_fd_sc_hd__buf_1
X_11497_ _05553_ net1815 _06432_ VGND VGND VPWR VPWR _06466_ sky130_fd_sc_hd__mux2_1
X_16024_ _02797_ _03502_ _03503_ _03504_ _02807_ VGND VGND VPWR VPWR _03505_ sky130_fd_sc_hd__a221o_1
X_13236_ CPU.registerFile\[15\]\[9\] _07402_ _07500_ CPU.registerFile\[11\]\[9\] _07327_
+ VGND VGND VPWR VPWR _07670_ sky130_fd_sc_hd__o221a_1
X_10448_ net1365 _05850_ _05851_ _05863_ VGND VGND VPWR VPWR _05864_ sky130_fd_sc_hd__a211o_1
Xclkbuf_1_1__f__02662_ clknet_0__02662_ VGND VGND VPWR VPWR clknet_1_1__leaf__02662_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_21_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__02693_ _02693_ VGND VGND VPWR VPWR clknet_0__02693_ sky130_fd_sc_hd__clkbuf_16
X_13167_ CPU.registerFile\[18\]\[8\] CPU.registerFile\[22\]\[8\] _07457_ VGND VGND
+ VPWR VPWR _07602_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10379_ _05811_ VGND VGND VPWR VPWR _02239_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__07220_ _07220_ VGND VGND VPWR VPWR clknet_0__07220_ sky130_fd_sc_hd__clkbuf_16
X_12118_ _06831_ VGND VGND VPWR VPWR _01516_ sky130_fd_sc_hd__clkbuf_1
X_17975_ net1163 _02259_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_13098_ CPU.registerFile\[23\]\[6\] _07236_ _07239_ CPU.registerFile\[19\]\[6\] _07534_
+ VGND VGND VPWR VPWR _07535_ sky130_fd_sc_hd__o221a_1
XFILLER_0_46_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12049_ _04982_ net2135 _06794_ VGND VGND VPWR VPWR _06795_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16857_ net1825 per_uart.rx_data\[7\] _04139_ VGND VGND VPWR VPWR _04147_ sky130_fd_sc_hd__mux2_1
X_15808_ _02948_ _03292_ _03295_ VGND VGND VPWR VPWR _03296_ sky130_fd_sc_hd__or3_2
X_16788_ _04050_ _04097_ _04098_ _04099_ VGND VGND VPWR VPWR _04100_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15739_ _02822_ VGND VGND VPWR VPWR _03228_ sky130_fd_sc_hd__buf_4
X_09260_ mapped_spi_ram.rcv_data\[13\] _04689_ _04691_ mapped_spi_flash.rcv_data\[13\]
+ VGND VGND VPWR VPWR _04970_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_158_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09191_ CPU.PC\[18\] _04836_ VGND VGND VPWR VPWR _04903_ sky130_fd_sc_hd__or2_1
X_17409_ net598 _01697_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_310 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__08467_ _08467_ VGND VGND VPWR VPWR clknet_0__08467_ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f__08367_ clknet_0__08367_ VGND VGND VPWR VPWR clknet_1_1__leaf__08367_
+ sky130_fd_sc_hd__clkbuf_16
X_08975_ CPU.Bimm\[10\] _04498_ _04687_ CPU.cycles\[30\] _04693_ VGND VGND VPWR VPWR
+ _04694_ sky130_fd_sc_hd__a221o_1
X_14249__421 clknet_1_0__leaf__08435_ VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__02751_ clknet_0__02751_ VGND VGND VPWR VPWR clknet_1_0__leaf__02751_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__02682_ clknet_0__02682_ VGND VGND VPWR VPWR clknet_1_0__leaf__02682_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_84_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09527_ _04888_ _05224_ VGND VGND VPWR VPWR _05225_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09458_ _04401_ _04430_ VGND VGND VPWR VPWR _05159_ sky130_fd_sc_hd__or2_1
X_09389_ _05092_ VGND VGND VPWR VPWR _05093_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_81_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14557__675 clknet_1_1__leaf__02671_ VGND VGND VPWR VPWR net707 sky130_fd_sc_hd__inv_2
X_11420_ _06425_ VGND VGND VPWR VPWR _01812_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11351_ _06388_ VGND VGND VPWR VPWR _01844_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10302_ _05770_ VGND VGND VPWR VPWR _02290_ sky130_fd_sc_hd__clkbuf_1
X_11282_ CPU.registerFile\[9\]\[6\] _05723_ _06346_ VGND VGND VPWR VPWR _06352_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13021_ CPU.registerFile\[23\]\[4\] _07362_ _07363_ CPU.registerFile\[19\]\[4\] _07459_
+ VGND VGND VPWR VPWR _07460_ sky130_fd_sc_hd__o221a_2
X_10233_ net2404 _05731_ _05713_ VGND VGND VPWR VPWR _05732_ sky130_fd_sc_hd__mux2_1
X_10164_ _04797_ VGND VGND VPWR VPWR _05685_ sky130_fd_sc_hd__clkbuf_4
X_15016__1089 clknet_1_1__leaf__02716_ VGND VGND VPWR VPWR net1121 sky130_fd_sc_hd__inv_2
X_17760_ net949 _02044_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_10095_ net1920 _04982_ _05644_ VGND VGND VPWR VPWR _05645_ sky130_fd_sc_hd__mux2_1
X_16711_ _05226_ _08454_ _05288_ VGND VGND VPWR VPWR _04035_ sky130_fd_sc_hd__and3b_1
X_13923_ CPU.registerFile\[16\]\[31\] CPU.registerFile\[20\]\[31\] _07648_ VGND VGND
+ VPWR VPWR _08335_ sky130_fd_sc_hd__mux2_1
X_14722__823 clknet_1_0__leaf__02688_ VGND VGND VPWR VPWR net855 sky130_fd_sc_hd__inv_2
X_17691_ net880 _01979_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_13854_ CPU.registerFile\[3\]\[29\] _07804_ _07987_ VGND VGND VPWR VPWR _08268_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12805_ CPU.registerFile\[21\]\[0\] _07244_ _07239_ CPU.registerFile\[17\]\[0\] _07247_
+ VGND VGND VPWR VPWR _07248_ sky130_fd_sc_hd__o221a_1
X_13785_ _07475_ _08200_ _08201_ VGND VGND VPWR VPWR _08202_ sky130_fd_sc_hd__o21a_1
X_10997_ _06200_ VGND VGND VPWR VPWR _02010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15524_ _08396_ VGND VGND VPWR VPWR _03019_ sky130_fd_sc_hd__buf_4
X_18312_ clknet_leaf_16_clk _02592_ VGND VGND VPWR VPWR CPU.PC\[12\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_128_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12736_ _07213_ net1575 _07205_ VGND VGND VPWR VPWR _07214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16596__67 clknet_1_1__leaf__03970_ VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__inv_2
XFILLER_0_57_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_106_Left_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18243_ net84 _02523_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15455_ _05050_ _02950_ _02951_ VGND VGND VPWR VPWR _02952_ sky130_fd_sc_hd__o21a_1
XFILLER_0_26_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12667_ CPU.cycles\[19\] _07158_ net1379 VGND VGND VPWR VPWR _07161_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18174_ net205 _02454_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_11618_ _06490_ _06547_ _06548_ _05942_ VGND VGND VPWR VPWR _01733_ sky130_fd_sc_hd__o31a_1
XFILLER_0_5_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15386_ _02882_ _02883_ _08400_ VGND VGND VPWR VPWR _02884_ sky130_fd_sc_hd__mux2_1
X_12598_ net1498 _07121_ _07122_ _07123_ _05815_ VGND VGND VPWR VPWR _00001_ sky130_fd_sc_hd__a221o_1
XFILLER_0_80_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17125_ clknet_leaf_20_clk _00028_ VGND VGND VPWR VPWR CPU.cycles\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11549_ _06501_ _04601_ VGND VGND VPWR VPWR _06502_ sky130_fd_sc_hd__nor2_1
Xhold507 CPU.registerFile\[4\]\[30\] VGND VGND VPWR VPWR net1748 sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 CPU.registerFile\[15\]\[25\] VGND VGND VPWR VPWR net1759 sky130_fd_sc_hd__dlygate4sd3_1
X_17056_ net314 _01378_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[18\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__02714_ clknet_0__02714_ VGND VGND VPWR VPWR clknet_1_1__leaf__02714_
+ sky130_fd_sc_hd__clkbuf_16
Xhold529 CPU.registerFile\[16\]\[0\] VGND VGND VPWR VPWR net1770 sky130_fd_sc_hd__dlygate4sd3_1
X_14268_ _08446_ _04674_ _04482_ _04481_ VGND VGND VPWR VPWR _08447_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_0_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16007_ CPU.registerFile\[31\]\[17\] _03072_ VGND VGND VPWR VPWR _03489_ sky130_fd_sc_hd__or2_1
X_13219_ _07272_ VGND VGND VPWR VPWR _07653_ sky130_fd_sc_hd__buf_6
Xclkbuf_0__02745_ _02745_ VGND VGND VPWR VPWR clknet_0__02745_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_122_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_115_Left_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__02676_ _02676_ VGND VGND VPWR VPWR clknet_0__02676_ sky130_fd_sc_hd__clkbuf_16
Xhold1207 CPU.rs2\[9\] VGND VGND VPWR VPWR net2448 sky130_fd_sc_hd__dlygate4sd3_1
X_08760_ _04479_ _04221_ VGND VGND VPWR VPWR _04480_ sky130_fd_sc_hd__nor2_1
Xhold1218 CPU.registerFile\[20\]\[20\] VGND VGND VPWR VPWR net2459 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17958_ net1146 _02242_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[3\] sky130_fd_sc_hd__dfxtp_1
Xhold1229 CPU.aluReg\[20\] VGND VGND VPWR VPWR net2470 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16909_ net1656 _04180_ _04183_ _04176_ VGND VGND VPWR VPWR _02638_ sky130_fd_sc_hd__o211a_1
X_08691_ _04297_ _04299_ _04290_ VGND VGND VPWR VPWR _04411_ sky130_fd_sc_hd__a21o_1
X_17889_ net1078 _02173_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_49_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_124_Left_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15033__1104 clknet_1_1__leaf__02718_ VGND VGND VPWR VPWR net1136 sky130_fd_sc_hd__inv_2
X_09312_ _04340_ _04699_ _04808_ CPU.aluReg\[19\] _05019_ VGND VGND VPWR VPWR _05020_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_87_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_815 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09243_ _04929_ _04953_ VGND VGND VPWR VPWR _04954_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09174_ CPU.Bimm\[8\] _04820_ CPU.PC\[8\] VGND VGND VPWR VPWR _04886_ sky130_fd_sc_hd__a21o_1
XFILLER_0_113_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15048__1115 clknet_1_0__leaf__02721_ VGND VGND VPWR VPWR net1147 sky130_fd_sc_hd__inv_2
XFILLER_0_32_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_133_Left_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08958_ CPU.Jimm\[14\] _04484_ VGND VGND VPWR VPWR _04677_ sky130_fd_sc_hd__nor2_1
X_08889_ _04564_ _04568_ _04569_ VGND VGND VPWR VPWR _04609_ sky130_fd_sc_hd__and3_1
X_10920_ net1675 _05702_ _06154_ VGND VGND VPWR VPWR _06160_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10851_ net2286 _05702_ _06117_ VGND VGND VPWR VPWR _06123_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__02665_ clknet_0__02665_ VGND VGND VPWR VPWR clknet_1_0__leaf__02665_
+ sky130_fd_sc_hd__clkbuf_16
X_15140__1169 clknet_1_0__leaf__02744_ VGND VGND VPWR VPWR net1201 sky130_fd_sc_hd__inv_2
X_13570_ CPU.registerFile\[18\]\[20\] CPU.registerFile\[22\]\[20\] _07457_ VGND VGND
+ VPWR VPWR _07993_ sky130_fd_sc_hd__mux2_1
X_10782_ _06086_ VGND VGND VPWR VPWR _02111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12521_ net1780 _05733_ _07048_ VGND VGND VPWR VPWR _07082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12452_ _07045_ VGND VGND VPWR VPWR _01362_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_10_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11403_ _06416_ VGND VGND VPWR VPWR _01820_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_97_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12383_ _05402_ net1937 _06999_ VGND VGND VPWR VPWR _07009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14122_ _08390_ VGND VGND VPWR VPWR _01469_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11334_ _06379_ VGND VGND VPWR VPWR _01852_ sky130_fd_sc_hd__clkbuf_1
X_11265_ CPU.registerFile\[9\]\[14\] _05706_ _06335_ VGND VGND VPWR VPWR _06343_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13004_ _07273_ _07442_ _07443_ VGND VGND VPWR VPWR _07444_ sky130_fd_sc_hd__o21a_1
X_10216_ _05720_ VGND VGND VPWR VPWR _02326_ sky130_fd_sc_hd__clkbuf_1
X_11196_ _06306_ VGND VGND VPWR VPWR _01917_ sky130_fd_sc_hd__clkbuf_1
X_17812_ net1001 _02096_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_10147_ net2093 _05673_ _05671_ VGND VGND VPWR VPWR _05674_ sky130_fd_sc_hd__mux2_1
X_14310__452 clknet_1_1__leaf__08464_ VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_128_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17743_ net932 _02027_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_10078_ net1621 _04714_ _05633_ VGND VGND VPWR VPWR _05636_ sky130_fd_sc_hd__mux2_1
X_13906_ CPU.registerFile\[29\]\[30\] _07502_ _07348_ CPU.registerFile\[25\]\[30\]
+ _07300_ VGND VGND VPWR VPWR _08319_ sky130_fd_sc_hd__o221a_1
X_17674_ net863 _01962_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[28\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_18_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13837_ _07273_ _08250_ _08251_ VGND VGND VPWR VPWR _08252_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_141_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13768_ CPU.registerFile\[16\]\[26\] CPU.registerFile\[20\]\[26\] _07258_ VGND VGND
+ VPWR VPWR _08185_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12719_ per_uart.uart0.tx_bitcount\[3\] per_uart.uart0.tx_bitcount\[2\] per_uart.uart0.tx_bitcount\[1\]
+ per_uart.uart0.tx_bitcount\[0\] VGND VGND VPWR VPWR _07201_ sky130_fd_sc_hd__or4_1
X_15507_ CPU.registerFile\[15\]\[4\] _02826_ _02770_ _03001_ VGND VGND VPWR VPWR _03002_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16487_ _03015_ _03952_ _03953_ _03954_ _02930_ VGND VGND VPWR VPWR _03955_ sky130_fd_sc_hd__a221o_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_13699_ CPU.registerFile\[1\]\[24\] _07387_ _08117_ _07379_ VGND VGND VPWR VPWR _08118_
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_44_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18226_ net67 _02506_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_15438_ _02934_ VGND VGND VPWR VPWR _02935_ sky130_fd_sc_hd__buf_2
XFILLER_0_143_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15369_ _02814_ VGND VGND VPWR VPWR _02867_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_14_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18157_ clknet_leaf_26_clk _02437_ VGND VGND VPWR VPWR CPU.aluIn1\[23\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_53_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold304 CPU.registerFile\[5\]\[1\] VGND VGND VPWR VPWR net1545 sky130_fd_sc_hd__dlygate4sd3_1
X_17108_ clknet_leaf_23_clk _00041_ VGND VGND VPWR VPWR CPU.cycles\[4\] sky130_fd_sc_hd__dfxtp_1
X_18088_ net151 _02368_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[18\] sky130_fd_sc_hd__dfxtp_1
Xhold315 CPU.registerFile\[18\]\[4\] VGND VGND VPWR VPWR net1556 sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 CPU.registerFile\[5\]\[12\] VGND VGND VPWR VPWR net1567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 CPU.registerFile\[28\]\[11\] VGND VGND VPWR VPWR net1578 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 CPU.registerFile\[6\]\[0\] VGND VGND VPWR VPWR net1589 sky130_fd_sc_hd__dlygate4sd3_1
X_09930_ _05447_ VGND VGND VPWR VPWR _05555_ sky130_fd_sc_hd__buf_4
X_17039_ net297 _01361_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold359 CPU.registerFile\[16\]\[1\] VGND VGND VPWR VPWR net1600 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09861_ _05508_ VGND VGND VPWR VPWR _02501_ sky130_fd_sc_hd__clkbuf_1
X_08812_ _04531_ _04530_ VGND VGND VPWR VPWR _04532_ sky130_fd_sc_hd__nand2_2
Xclkbuf_0__02659_ _02659_ VGND VGND VPWR VPWR clknet_0__02659_ sky130_fd_sc_hd__clkbuf_16
Xhold1004 CPU.registerFile\[20\]\[3\] VGND VGND VPWR VPWR net2245 sky130_fd_sc_hd__dlygate4sd3_1
X_09792_ net2535 _05046_ _05463_ VGND VGND VPWR VPWR _05467_ sky130_fd_sc_hd__mux2_1
Xhold1015 CPU.registerFile\[17\]\[14\] VGND VGND VPWR VPWR net2256 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1026 CPU.registerFile\[18\]\[17\] VGND VGND VPWR VPWR net2267 sky130_fd_sc_hd__dlygate4sd3_1
X_08743_ _04462_ _04382_ _04350_ VGND VGND VPWR VPWR _04463_ sky130_fd_sc_hd__o21bai_1
Xhold1037 CPU.registerFile\[17\]\[15\] VGND VGND VPWR VPWR net2278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1048 CPU.PC\[8\] VGND VGND VPWR VPWR net2289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 CPU.registerFile\[10\]\[2\] VGND VGND VPWR VPWR net2300 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08674_ _04393_ _04257_ VGND VGND VPWR VPWR _04394_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16575__48 clknet_1_0__leaf__03968_ VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__inv_2
X_09226_ _04936_ VGND VGND VPWR VPWR _04937_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15015__1088 clknet_1_1__leaf__02716_ VGND VGND VPWR VPWR net1120 sky130_fd_sc_hd__inv_2
XFILLER_0_134_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09157_ CPU.PC\[3\] _04868_ VGND VGND VPWR VPWR _04869_ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_141_Left_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09088_ _04670_ VGND VGND VPWR VPWR _04800_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold860 CPU.registerFile\[17\]\[22\] VGND VGND VPWR VPWR net2101 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold871 CPU.registerFile\[19\]\[9\] VGND VGND VPWR VPWR net2112 sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 CPU.registerFile\[29\]\[17\] VGND VGND VPWR VPWR net2123 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14669__776 clknet_1_0__leaf__02682_ VGND VGND VPWR VPWR net808 sky130_fd_sc_hd__inv_2
X_11050_ CPU.registerFile\[7\]\[19\] _05696_ _06226_ VGND VGND VPWR VPWR _06229_ sky130_fd_sc_hd__mux2_1
Xhold893 CPU.registerFile\[28\]\[24\] VGND VGND VPWR VPWR net2134 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10001_ _05593_ VGND VGND VPWR VPWR _02446_ sky130_fd_sc_hd__clkbuf_1
X_14740_ clknet_1_0__leaf__02686_ VGND VGND VPWR VPWR _02690_ sky130_fd_sc_hd__buf_1
X_11952_ CPU.registerFile\[11\]\[2\] _05731_ _06733_ VGND VGND VPWR VPWR _06743_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10903_ net1727 _05685_ _06143_ VGND VGND VPWR VPWR _06151_ sky130_fd_sc_hd__mux2_1
X_11883_ _06706_ VGND VGND VPWR VPWR _01627_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__02717_ clknet_0__02717_ VGND VGND VPWR VPWR clknet_1_0__leaf__02717_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_123_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16410_ CPU.registerFile\[10\]\[29\] _02928_ _02910_ VGND VGND VPWR VPWR _03880_
+ sky130_fd_sc_hd__o21a_1
X_13622_ CPU.registerFile\[2\]\[21\] _07388_ VGND VGND VPWR VPWR _08044_ sky130_fd_sc_hd__or2_1
XFILLER_0_157_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10834_ net1658 _05685_ _06106_ VGND VGND VPWR VPWR _06114_ sky130_fd_sc_hd__mux2_1
X_17390_ net579 _01678_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16341_ CPU.registerFile\[16\]\[27\] CPU.registerFile\[20\]\[27\] _02777_ VGND VGND
+ VPWR VPWR _03813_ sky130_fd_sc_hd__mux2_1
X_14834__924 clknet_1_1__leaf__02699_ VGND VGND VPWR VPWR net956 sky130_fd_sc_hd__inv_2
X_13553_ CPU.registerFile\[28\]\[19\] CPU.registerFile\[24\]\[19\] _07399_ VGND VGND
+ VPWR VPWR _07977_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10765_ _06077_ VGND VGND VPWR VPWR _02119_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12504_ _07073_ VGND VGND VPWR VPWR _01338_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16272_ _02767_ _03741_ _03745_ _05361_ VGND VGND VPWR VPWR _03746_ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13484_ CPU.registerFile\[23\]\[17\] _07325_ _07500_ CPU.registerFile\[19\]\[17\]
+ _07327_ VGND VGND VPWR VPWR _07910_ sky130_fd_sc_hd__o221a_1
XFILLER_0_82_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10696_ _05503_ net2445 _06034_ VGND VGND VPWR VPWR _06041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18011_ net1184 _02291_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12435_ _05209_ net2017 _07035_ VGND VGND VPWR VPWR _07037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_391 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12366_ _07000_ VGND VGND VPWR VPWR _01403_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_136_Right_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14105_ _04292_ _05340_ _00000_ VGND VGND VPWR VPWR _08381_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11317_ _06370_ VGND VGND VPWR VPWR _01860_ sky130_fd_sc_hd__clkbuf_1
X_15085_ _02729_ VGND VGND VPWR VPWR _02272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12297_ CPU.aluReg\[6\] CPU.aluReg\[4\] _06939_ VGND VGND VPWR VPWR _06958_ sky130_fd_sc_hd__mux2_1
X_15032__1103 clknet_1_1__leaf__02718_ VGND VGND VPWR VPWR net1135 sky130_fd_sc_hd__inv_2
X_11248_ net2320 _05689_ _06324_ VGND VGND VPWR VPWR _06334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14880__966 clknet_1_0__leaf__02703_ VGND VGND VPWR VPWR net998 sky130_fd_sc_hd__inv_2
X_11179_ _06297_ VGND VGND VPWR VPWR _01925_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_143_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15987_ _03465_ _03468_ _08401_ VGND VGND VPWR VPWR _03469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15047__1114 clknet_1_1__leaf__02721_ VGND VGND VPWR VPWR net1146 sky130_fd_sc_hd__inv_2
X_17726_ net915 _02010_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17657_ net846 _01945_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16608_ _03978_ VGND VGND VPWR VPWR _03979_ sky130_fd_sc_hd__buf_2
X_17588_ net777 _01876_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_158_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09011_ _04362_ _04489_ _04727_ _04679_ VGND VGND VPWR VPWR _04728_ sky130_fd_sc_hd__a22o_1
X_18209_ net50 _02489_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_154_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold101 _01327_ VGND VGND VPWR VPWR net1342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 _02276_ VGND VGND VPWR VPWR net1353 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 _02271_ VGND VGND VPWR VPWR net1364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_103_Right_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold134 mapped_spi_ram.cmd_addr\[11\] VGND VGND VPWR VPWR net1375 sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 mapped_spi_ram.cmd_addr\[14\] VGND VGND VPWR VPWR net1386 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 mapped_spi_flash.cmd_addr\[12\] VGND VGND VPWR VPWR net1397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 _01725_ VGND VGND VPWR VPWR net1408 sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ _05543_ net2531 _05533_ VGND VGND VPWR VPWR _05544_ sky130_fd_sc_hd__mux2_1
Xhold178 CPU.cycles\[2\] VGND VGND VPWR VPWR net1419 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold189 mapped_spi_flash.snd_bitcount\[4\] VGND VGND VPWR VPWR net1430 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09844_ _04730_ VGND VGND VPWR VPWR _05497_ sky130_fd_sc_hd__clkbuf_4
X_09775_ net1828 _04762_ _05452_ VGND VGND VPWR VPWR _05458_ sky130_fd_sc_hd__mux2_1
X_15218__129 clknet_1_0__leaf__02752_ VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__inv_2
X_08726_ _04388_ _04443_ _04445_ VGND VGND VPWR VPWR _04446_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_1_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ CPU.aluIn1\[29\] VGND VGND VPWR VPWR _04377_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08588_ CPU.aluIn1\[4\] _04284_ VGND VGND VPWR VPWR _04308_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10550_ _05886_ _05946_ _05947_ net1418 VGND VGND VPWR VPWR _05948_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09209_ CPU.PC\[10\] CPU.PC\[9\] _04920_ VGND VGND VPWR VPWR _04921_ sky130_fd_sc_hd__and3_1
XFILLER_0_106_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10481_ net1397 _05849_ _05891_ _05885_ VGND VGND VPWR VPWR _02216_ sky130_fd_sc_hd__o211a_1
X_12220_ _06899_ VGND VGND VPWR VPWR _01448_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_20_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12151_ _06848_ VGND VGND VPWR VPWR _01500_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11102_ net1740 _05679_ _06252_ VGND VGND VPWR VPWR _06257_ sky130_fd_sc_hd__mux2_1
X_12082_ _05333_ net2071 _06805_ VGND VGND VPWR VPWR _06812_ sky130_fd_sc_hd__mux2_1
Xhold690 CPU.registerFile\[20\]\[13\] VGND VGND VPWR VPWR net1931 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11033_ net1617 _05679_ _06215_ VGND VGND VPWR VPWR _06220_ sky130_fd_sc_hd__mux2_1
X_15910_ _02926_ _03393_ _03394_ VGND VGND VPWR VPWR _03395_ sky130_fd_sc_hd__o21a_1
X_16890_ net1839 _04168_ _04170_ _03632_ VGND VGND VPWR VPWR _02632_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_125_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15841_ CPU.registerFile\[18\]\[12\] _02832_ _02835_ CPU.registerFile\[19\]\[12\]
+ _03074_ VGND VGND VPWR VPWR _03328_ sky130_fd_sc_hd__o221a_1
X_12984_ _07397_ _07410_ _07423_ _07424_ VGND VGND VPWR VPWR _07425_ sky130_fd_sc_hd__a31o_1
X_15772_ CPU.registerFile\[30\]\[10\] _05050_ _02923_ _03260_ VGND VGND VPWR VPWR
+ _03261_ sky130_fd_sc_hd__o211a_1
X_17511_ net700 _01799_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_11935_ _06734_ VGND VGND VPWR VPWR _01603_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_748 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17442_ net631 _01730_ VGND VGND VPWR VPWR mapped_spi_ram.snd_bitcount\[3\] sky130_fd_sc_hd__dfxtp_1
X_11866_ net2381 _05712_ _06697_ VGND VGND VPWR VPWR _06698_ sky130_fd_sc_hd__mux2_1
X_16539__15 clknet_1_0__leaf__03965_ VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__inv_2
X_14422__553 clknet_1_0__leaf__02658_ VGND VGND VPWR VPWR net585 sky130_fd_sc_hd__inv_2
X_13605_ _07370_ _08026_ VGND VGND VPWR VPWR _08027_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10817_ _06104_ VGND VGND VPWR VPWR _02094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17373_ net562 _01661_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11797_ _06638_ VGND VGND VPWR VPWR _06661_ sky130_fd_sc_hd__buf_4
XFILLER_0_131_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16324_ CPU.registerFile\[8\]\[27\] CPU.registerFile\[12\]\[27\] _02852_ VGND VGND
+ VPWR VPWR _03796_ sky130_fd_sc_hd__mux2_1
X_13536_ _07288_ _07959_ VGND VGND VPWR VPWR _07960_ sky130_fd_sc_hd__or2_1
X_10748_ _05555_ net1653 _06033_ VGND VGND VPWR VPWR _06068_ sky130_fd_sc_hd__mux2_1
X_16554__29 clknet_1_1__leaf__03966_ VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__inv_2
XFILLER_0_125_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16255_ _08407_ _03706_ _03715_ _03729_ _07424_ VGND VGND VPWR VPWR _03730_ sky130_fd_sc_hd__a311o_1
X_13467_ CPU.rs2\[16\] _07705_ _07878_ _07893_ _07737_ VGND VGND VPWR VPWR _01311_
+ sky130_fd_sc_hd__o221a_1
X_10679_ net1314 _06010_ VGND VGND VPWR VPWR _06031_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_136_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12418_ net1245 net1861 _07024_ VGND VGND VPWR VPWR _07028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16186_ _03659_ _03660_ _03662_ _02812_ VGND VGND VPWR VPWR _03663_ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13398_ _07291_ _07826_ VGND VGND VPWR VPWR _07827_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12349_ _06991_ VGND VGND VPWR VPWR _01411_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15014__1087 clknet_1_1__leaf__02716_ VGND VGND VPWR VPWR net1119 sky130_fd_sc_hd__inv_2
XFILLER_0_65_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09560_ _04884_ _04861_ VGND VGND VPWR VPWR _05256_ sky130_fd_sc_hd__or2b_1
X_08511_ CPU.rs2\[26\] _04201_ _04206_ VGND VGND VPWR VPWR _04231_ sky130_fd_sc_hd__a21o_1
X_14505__628 clknet_1_1__leaf__02666_ VGND VGND VPWR VPWR net660 sky130_fd_sc_hd__inv_2
X_17709_ net898 _01997_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_09491_ _05190_ VGND VGND VPWR VPWR _02561_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14243__416 clknet_1_0__leaf__08434_ VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__inv_2
XFILLER_0_147_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_156_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14397__530 clknet_1_0__leaf__02656_ VGND VGND VPWR VPWR net562 sky130_fd_sc_hd__inv_2
XFILLER_0_73_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14863__950 clknet_1_0__leaf__02702_ VGND VGND VPWR VPWR net982 sky130_fd_sc_hd__inv_2
XFILLER_0_10_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09827_ net2024 _05426_ _05451_ VGND VGND VPWR VPWR _05485_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09758_ _04492_ _05438_ _05446_ VGND VGND VPWR VPWR _05447_ sky130_fd_sc_hd__a21o_2
X_08709_ _04403_ _04427_ _04428_ VGND VGND VPWR VPWR _04429_ sky130_fd_sc_hd__o21a_1
XFILLER_0_69_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09689_ _05380_ VGND VGND VPWR VPWR _05381_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_87_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11720_ net1473 _06603_ _06614_ _06607_ VGND VGND VPWR VPWR _01697_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_120_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ _06574_ VGND VGND VPWR VPWR _06575_ sky130_fd_sc_hd__buf_2
X_15031__1102 clknet_1_1__leaf__02718_ VGND VGND VPWR VPWR net1134 sky130_fd_sc_hd__inv_2
XFILLER_0_36_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10602_ mapped_spi_flash.rcv_data\[21\] _05981_ VGND VGND VPWR VPWR _05984_ sky130_fd_sc_hd__or2_1
X_11582_ net1386 _06524_ _06516_ _06526_ VGND VGND VPWR VPWR _01747_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13321_ _07232_ _07744_ _07751_ VGND VGND VPWR VPWR _07752_ sky130_fd_sc_hd__a21o_1
XFILLER_0_92_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10533_ net1442 _05887_ _05856_ _05934_ VGND VGND VPWR VPWR _05935_ sky130_fd_sc_hd__a211o_1
XFILLER_0_51_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16040_ _03517_ _03518_ _03520_ _02812_ VGND VGND VPWR VPWR _03521_ sky130_fd_sc_hd__o22a_2
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13252_ CPU.registerFile\[21\]\[10\] _07403_ _07619_ CPU.registerFile\[17\]\[10\]
+ _07250_ VGND VGND VPWR VPWR _07685_ sky130_fd_sc_hd__o221a_1
X_10464_ _04629_ _05868_ _05875_ _05876_ VGND VGND VPWR VPWR _05877_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_118_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15046__1113 clknet_1_1__leaf__02721_ VGND VGND VPWR VPWR net1145 sky130_fd_sc_hd__inv_2
XFILLER_0_20_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12203_ CPU.aluReg\[28\] CPU.aluReg\[26\] _06871_ VGND VGND VPWR VPWR _06886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13183_ _07238_ VGND VGND VPWR VPWR _07618_ sky130_fd_sc_hd__clkbuf_8
X_10395_ _05824_ VGND VGND VPWR VPWR _05825_ sky130_fd_sc_hd__buf_2
XFILLER_0_103_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12134_ _06839_ VGND VGND VPWR VPWR _01508_ sky130_fd_sc_hd__clkbuf_1
X_17991_ clknet_leaf_10_clk _02275_ VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_16942_ net237 _01268_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_12065_ _05150_ net2169 _06794_ VGND VGND VPWR VPWR _06803_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11016_ _06210_ VGND VGND VPWR VPWR _02001_ sky130_fd_sc_hd__clkbuf_1
X_16873_ _04156_ _04157_ _04158_ VGND VGND VPWR VPWR _04159_ sky130_fd_sc_hd__o21a_1
XFILLER_0_126_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15824_ _02911_ _03308_ _03310_ _02794_ VGND VGND VPWR VPWR _03311_ sky130_fd_sc_hd__a211o_1
X_15755_ CPU.registerFile\[10\]\[10\] _02816_ _02910_ VGND VGND VPWR VPWR _03244_
+ sky130_fd_sc_hd__o21a_1
X_12967_ CPU.registerFile\[28\]\[2\] CPU.registerFile\[24\]\[2\] _07399_ VGND VGND
+ VPWR VPWR _07408_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14706_ clknet_1_0__leaf__07222_ VGND VGND VPWR VPWR _02686_ sky130_fd_sc_hd__buf_1
X_11918_ _06725_ VGND VGND VPWR VPWR _01611_ sky130_fd_sc_hd__clkbuf_1
X_15686_ CPU.registerFile\[5\]\[8\] CPU.registerFile\[4\]\[8\] _02805_ VGND VGND VPWR
+ VPWR _03177_ sky130_fd_sc_hd__mux2_1
X_12898_ CPU.registerFile\[8\]\[1\] CPU.registerFile\[12\]\[1\] _07339_ VGND VGND
+ VPWR VPWR _07340_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_360 _07291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_371 _05381_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_382 _05272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17425_ net614 net1436 VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_393 _07318_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11849_ CPU.registerFile\[10\]\[19\] _05696_ _06686_ VGND VGND VPWR VPWR _06689_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17356_ net545 _01644_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16307_ CPU.registerFile\[30\]\[26\] CPU.registerFile\[26\]\[26\] _02773_ VGND VGND
+ VPWR VPWR _03780_ sky130_fd_sc_hd__mux2_1
X_13519_ _07418_ _07942_ _07943_ VGND VGND VPWR VPWR _07944_ sky130_fd_sc_hd__o21a_1
X_17287_ net476 _01575_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_15247__155 clknet_1_0__leaf__02755_ VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__inv_2
Xclkload10 clknet_leaf_13_clk VGND VGND VPWR VPWR clkload10/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_151_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload21 clknet_leaf_5_clk VGND VGND VPWR VPWR clkload21/Y sky130_fd_sc_hd__clkinv_4
X_16238_ CPU.registerFile\[25\]\[24\] _03280_ _02940_ VGND VGND VPWR VPWR _03713_
+ sky130_fd_sc_hd__o21a_1
Xclkload32 clknet_1_0__leaf__02754_ VGND VGND VPWR VPWR clkload32/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload43 clknet_1_1__leaf__02724_ VGND VGND VPWR VPWR clkload43/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_2_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload54 clknet_1_1__leaf__02703_ VGND VGND VPWR VPWR clkload54/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload65 clknet_1_0__leaf__02675_ VGND VGND VPWR VPWR clkload65/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_51_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload76 clknet_1_1__leaf__02668_ VGND VGND VPWR VPWR clkload76/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_141_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload87 clknet_1_1__leaf__02657_ VGND VGND VPWR VPWR clkload87/Y sky130_fd_sc_hd__clkinvlp_4
X_16169_ CPU.registerFile\[29\]\[22\] _02926_ VGND VGND VPWR VPWR _03646_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload98 clknet_1_0__leaf__08431_ VGND VGND VPWR VPWR clkload98/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_54_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08991_ _04690_ VGND VGND VPWR VPWR _04709_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_54_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14585__700 clknet_1_0__leaf__02674_ VGND VGND VPWR VPWR net732 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_71_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09612_ net1777 _05306_ _05189_ VGND VGND VPWR VPWR _05307_ sky130_fd_sc_hd__mux2_1
X_09543_ CPU.PC\[8\] _04919_ VGND VGND VPWR VPWR _05240_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_69_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09474_ _04782_ _05172_ _05173_ _04681_ VGND VGND VPWR VPWR _05174_ sky130_fd_sc_hd__a22oi_2
XTAP_TAPCELL_ROW_102_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload4 clknet_leaf_24_clk VGND VGND VPWR VPWR clkload4/Y sky130_fd_sc_hd__inv_8
XFILLER_0_144_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_355 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10180_ _05026_ VGND VGND VPWR VPWR _05696_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13870_ CPU.registerFile\[8\]\[29\] CPU.registerFile\[12\]\[29\] _07339_ VGND VGND
+ VPWR VPWR _08284_ sky130_fd_sc_hd__mux2_1
X_12821_ CPU.registerFile\[6\]\[0\] _07263_ VGND VGND VPWR VPWR _07264_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15540_ _02903_ _03029_ _03034_ VGND VGND VPWR VPWR _03035_ sky130_fd_sc_hd__or3_1
XFILLER_0_29_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11703_ net2471 _06603_ _06605_ _06594_ VGND VGND VPWR VPWR _01705_ sky130_fd_sc_hd__o211a_1
X_15471_ _08397_ _02961_ _02963_ _02966_ VGND VGND VPWR VPWR _02967_ sky130_fd_sc_hd__o22a_1
X_12683_ CPU.cycles\[27\] _07168_ VGND VGND VPWR VPWR _07170_ sky130_fd_sc_hd__and2_1
X_17210_ net400 _01498_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_11634_ _06555_ VGND VGND VPWR VPWR _06562_ sky130_fd_sc_hd__inv_2
XFILLER_0_37_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18190_ net221 _02470_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17141_ net365 _01429_ VGND VGND VPWR VPWR CPU.aluReg\[5\] sky130_fd_sc_hd__dfxtp_1
X_11565_ net1358 _06499_ _06509_ _06513_ VGND VGND VPWR VPWR _06514_ sky130_fd_sc_hd__a211o_1
XFILLER_0_107_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13304_ _07397_ _07728_ _07735_ _07703_ VGND VGND VPWR VPWR _07736_ sky130_fd_sc_hd__a31o_1
X_15013__1086 clknet_1_1__leaf__02716_ VGND VGND VPWR VPWR net1118 sky130_fd_sc_hd__inv_2
X_17072_ net330 _01394_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_10516_ net1382 _05892_ _05921_ _05885_ VGND VGND VPWR VPWR _02211_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_133_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11496_ _06465_ VGND VGND VPWR VPWR _01776_ sky130_fd_sc_hd__clkbuf_1
X_14079__352 clknet_1_0__leaf__08368_ VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__inv_2
XFILLER_0_52_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14534__654 clknet_1_1__leaf__02669_ VGND VGND VPWR VPWR net686 sky130_fd_sc_hd__inv_2
XFILLER_0_134_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16023_ CPU.registerFile\[9\]\[18\] _02802_ _03125_ VGND VGND VPWR VPWR _03504_ sky130_fd_sc_hd__o21a_1
XFILLER_0_21_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13235_ CPU.registerFile\[14\]\[9\] CPU.registerFile\[10\]\[9\] _07492_ VGND VGND
+ VPWR VPWR _07669_ sky130_fd_sc_hd__mux2_1
X_10447_ _05852_ _04604_ VGND VGND VPWR VPWR _05863_ sky130_fd_sc_hd__nor2_1
Xclkbuf_1_1__f__02661_ clknet_0__02661_ VGND VGND VPWR VPWR clknet_1_1__leaf__02661_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_32_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13166_ CPU.mem_wdata\[7\] _07358_ _07586_ _07601_ _05844_ VGND VGND VPWR VPWR _01302_
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_0__02692_ _02692_ VGND VGND VPWR VPWR clknet_0__02692_ sky130_fd_sc_hd__clkbuf_16
X_10378_ _05555_ net2389 _05776_ VGND VGND VPWR VPWR _05811_ sky130_fd_sc_hd__mux2_1
X_12117_ _04982_ net2232 _06830_ VGND VGND VPWR VPWR _06831_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17974_ net1162 _02258_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_13097_ _05338_ _07533_ VGND VGND VPWR VPWR _07534_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12048_ _06782_ VGND VGND VPWR VPWR _06794_ sky130_fd_sc_hd__buf_4
XFILLER_0_137_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16856_ net1798 VGND VGND VPWR VPWR _02622_ sky130_fd_sc_hd__clkbuf_1
X_15807_ _03072_ _03293_ _03294_ VGND VGND VPWR VPWR _03295_ sky130_fd_sc_hd__o21a_1
X_16787_ _04914_ _04963_ _03990_ VGND VGND VPWR VPWR _04099_ sky130_fd_sc_hd__a21o_1
X_14580__696 clknet_1_0__leaf__02673_ VGND VGND VPWR VPWR net728 sky130_fd_sc_hd__inv_2
XFILLER_0_88_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15738_ _02821_ VGND VGND VPWR VPWR _03227_ sky130_fd_sc_hd__buf_4
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15669_ CPU.registerFile\[12\]\[8\] _03118_ VGND VGND VPWR VPWR _03160_ sky130_fd_sc_hd__or2_1
XANTENNA_190 _07841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17408_ net597 _01696_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_64_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09190_ _04841_ _04901_ _04839_ VGND VGND VPWR VPWR _04902_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_16_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14617__729 clknet_1_1__leaf__02677_ VGND VGND VPWR VPWR net761 sky130_fd_sc_hd__inv_2
XFILLER_0_145_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17339_ net528 _01627_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload110 clknet_1_1__leaf__07226_ VGND VGND VPWR VPWR clkload110/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__08435_ clknet_0__08435_ VGND VGND VPWR VPWR clknet_1_1__leaf__08435_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_140_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__08466_ _08466_ VGND VGND VPWR VPWR clknet_0__08466_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__08366_ clknet_0__08366_ VGND VGND VPWR VPWR clknet_1_1__leaf__08366_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08974_ _04216_ _04692_ _04655_ VGND VGND VPWR VPWR _04693_ sky130_fd_sc_hd__o21ba_1
X_15030__1101 clknet_1_0__leaf__02718_ VGND VGND VPWR VPWR net1133 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__02750_ clknet_0__02750_ VGND VGND VPWR VPWR clknet_1_0__leaf__02750_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15045__1112 clknet_1_0__leaf__02721_ VGND VGND VPWR VPWR net1144 sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__02681_ clknet_0__02681_ VGND VGND VPWR VPWR clknet_1_0__leaf__02681_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_84_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09526_ _04859_ _04887_ VGND VGND VPWR VPWR _05224_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09457_ _04433_ _04324_ VGND VGND VPWR VPWR _05158_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_913 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09388_ net15 VGND VGND VPWR VPWR _05092_ sky130_fd_sc_hd__buf_4
XFILLER_0_81_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11350_ _05543_ net2454 _06382_ VGND VGND VPWR VPWR _06388_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10301_ _05547_ net2314 _05762_ VGND VGND VPWR VPWR _05770_ sky130_fd_sc_hd__mux2_1
X_11281_ _06351_ VGND VGND VPWR VPWR _01877_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13020_ _07364_ _07458_ VGND VGND VPWR VPWR _07459_ sky130_fd_sc_hd__or2_1
X_10232_ _05401_ VGND VGND VPWR VPWR _05731_ sky130_fd_sc_hd__clkbuf_4
X_10163_ _05684_ VGND VGND VPWR VPWR _02343_ sky130_fd_sc_hd__clkbuf_1
X_10094_ _05632_ VGND VGND VPWR VPWR _05644_ sky130_fd_sc_hd__buf_4
X_16710_ _08436_ _08459_ _05225_ VGND VGND VPWR VPWR _04034_ sky130_fd_sc_hd__a21oi_1
X_13922_ CPU.registerFile\[23\]\[31\] _07282_ _08333_ VGND VGND VPWR VPWR _08334_
+ sky130_fd_sc_hd__o21ai_1
X_17690_ net879 _01978_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13853_ CPU.registerFile\[2\]\[29\] _07621_ VGND VGND VPWR VPWR _08267_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12804_ _07245_ _07246_ VGND VGND VPWR VPWR _07247_ sky130_fd_sc_hd__or2_1
X_10996_ net2518 _05710_ _06190_ VGND VGND VPWR VPWR _06200_ sky130_fd_sc_hd__mux2_1
X_13784_ CPU.registerFile\[15\]\[26\] _07325_ _07500_ CPU.registerFile\[11\]\[26\]
+ _07327_ VGND VGND VPWR VPWR _08201_ sky130_fd_sc_hd__o221a_1
XFILLER_0_69_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18311_ clknet_leaf_16_clk _02591_ VGND VGND VPWR VPWR CPU.PC\[11\] sky130_fd_sc_hd__dfxtp_1
X_15523_ _02796_ _03017_ VGND VGND VPWR VPWR _03018_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12735_ per_uart.d_in_uart\[2\] _07178_ _07203_ per_uart.uart0.txd_reg\[3\] VGND
+ VGND VPWR VPWR _07213_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18242_ net83 _02522_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12666_ CPU.cycles\[19\] CPU.cycles\[20\] _07158_ VGND VGND VPWR VPWR _07160_ sky130_fd_sc_hd__and3_1
X_15454_ CPU.registerFile\[16\]\[2\] _02832_ _02835_ CPU.registerFile\[17\]\[2\] _02940_
+ VGND VGND VPWR VPWR _02951_ sky130_fd_sc_hd__o221a_1
XFILLER_0_38_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11617_ CPU.mem_wdata\[0\] _06470_ _06487_ VGND VGND VPWR VPWR _06548_ sky130_fd_sc_hd__and3_1
X_18173_ net204 _02453_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_12597_ CPU.state\[1\] VGND VGND VPWR VPWR _07123_ sky130_fd_sc_hd__clkbuf_4
X_15385_ CPU.registerFile\[30\]\[1\] CPU.registerFile\[26\]\[1\] _02881_ VGND VGND
+ VPWR VPWR _02883_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17124_ clknet_leaf_17_clk _00027_ VGND VGND VPWR VPWR CPU.cycles\[20\] sky130_fd_sc_hd__dfxtp_1
X_11548_ _06493_ VGND VGND VPWR VPWR _06501_ sky130_fd_sc_hd__buf_2
Xhold508 CPU.registerFile\[30\]\[27\] VGND VGND VPWR VPWR net1749 sky130_fd_sc_hd__dlygate4sd3_1
X_14267_ _04704_ _04736_ _04751_ _08445_ VGND VGND VPWR VPWR _08446_ sky130_fd_sc_hd__or4_1
Xhold519 CPU.registerFile\[9\]\[30\] VGND VGND VPWR VPWR net1760 sky130_fd_sc_hd__dlygate4sd3_1
X_17055_ net313 _01377_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[17\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__02713_ clknet_0__02713_ VGND VGND VPWR VPWR clknet_1_1__leaf__02713_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11479_ _05535_ CPU.registerFile\[25\]\[10\] _06455_ VGND VGND VPWR VPWR _06457_
+ sky130_fd_sc_hd__mux2_1
X_16006_ CPU.registerFile\[25\]\[17\] CPU.registerFile\[29\]\[17\] _03254_ VGND VGND
+ VPWR VPWR _03488_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__02744_ _02744_ VGND VGND VPWR VPWR clknet_0__02744_ sky130_fd_sc_hd__clkbuf_16
X_13218_ CPU.registerFile\[19\]\[9\] _07383_ _07651_ VGND VGND VPWR VPWR _07652_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13149_ _07380_ _07579_ _07583_ _07584_ VGND VGND VPWR VPWR _07585_ sky130_fd_sc_hd__o211a_4
Xclkbuf_0__02675_ _02675_ VGND VGND VPWR VPWR clknet_0__02675_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1208 CPU.registerFile\[25\]\[9\] VGND VGND VPWR VPWR net2449 sky130_fd_sc_hd__dlygate4sd3_1
X_17957_ net1145 _02241_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[2\] sky130_fd_sc_hd__dfxtp_1
Xhold1219 CPU.registerFile\[7\]\[8\] VGND VGND VPWR VPWR net2460 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_146_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16908_ net1768 _04182_ VGND VGND VPWR VPWR _04183_ sky130_fd_sc_hd__or2_1
X_08690_ _04290_ _04409_ VGND VGND VPWR VPWR _04410_ sky130_fd_sc_hd__or2_1
X_17888_ net1077 net1396 VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[6\] sky130_fd_sc_hd__dfxtp_1
X_16839_ _04136_ _07203_ net1410 _06030_ VGND VGND VPWR VPWR _02615_ sky130_fd_sc_hd__a2bb2o_1
X_14697__801 clknet_1_1__leaf__02685_ VGND VGND VPWR VPWR net833 sky130_fd_sc_hd__inv_2
XFILLER_0_88_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_49_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09311_ _04447_ _04682_ VGND VGND VPWR VPWR _05019_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09242_ CPU.PC\[21\] _04928_ CPU.PC\[22\] VGND VGND VPWR VPWR _04953_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_907 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_778 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09173_ _04861_ _04883_ _04884_ VGND VGND VPWR VPWR _04885_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08957_ _04368_ _04675_ _04374_ VGND VGND VPWR VPWR _04676_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08888_ CPU.PC\[19\] _04586_ _04606_ _04607_ VGND VGND VPWR VPWR _04608_ sky130_fd_sc_hd__o2bb2a_1
X_15012__1085 clknet_1_0__leaf__02716_ VGND VGND VPWR VPWR net1117 sky130_fd_sc_hd__inv_2
X_14563__680 clknet_1_1__leaf__02672_ VGND VGND VPWR VPWR net712 sky130_fd_sc_hd__inv_2
X_10850_ _06122_ VGND VGND VPWR VPWR _02079_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__02664_ clknet_0__02664_ VGND VGND VPWR VPWR clknet_1_0__leaf__02664_
+ sky130_fd_sc_hd__clkbuf_16
X_09509_ CPU.cycles\[10\] _04687_ _05193_ _05207_ VGND VGND VPWR VPWR _05208_ sky130_fd_sc_hd__a211o_4
X_10781_ _05520_ net2172 _06081_ VGND VGND VPWR VPWR _06086_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12520_ _07081_ VGND VGND VPWR VPWR _01330_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_117_Right_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12451_ _05402_ net2283 _07035_ VGND VGND VPWR VPWR _07045_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_10_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11402_ _05526_ net2053 _06408_ VGND VGND VPWR VPWR _06416_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12382_ _07008_ VGND VGND VPWR VPWR _01395_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_97_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_90 _05305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14121_ _04665_ _08389_ _08387_ VGND VGND VPWR VPWR _08390_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11333_ _05526_ net2513 _06371_ VGND VGND VPWR VPWR _06379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11264_ _06342_ VGND VGND VPWR VPWR _01885_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13003_ CPU.registerFile\[15\]\[3\] _07276_ _07277_ CPU.registerFile\[11\]\[3\] _07278_
+ VGND VGND VPWR VPWR _07443_ sky130_fd_sc_hd__o221a_1
X_10215_ net2234 _05719_ _05713_ VGND VGND VPWR VPWR _05720_ sky130_fd_sc_hd__mux2_1
X_11195_ _05524_ net1643 _06299_ VGND VGND VPWR VPWR _06306_ sky130_fd_sc_hd__mux2_1
X_17811_ net1000 _02095_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_10146_ _04695_ VGND VGND VPWR VPWR _05673_ sky130_fd_sc_hd__buf_2
X_14646__755 clknet_1_1__leaf__02680_ VGND VGND VPWR VPWR net787 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_128_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17742_ net931 _02026_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_10077_ _05635_ VGND VGND VPWR VPWR _02380_ sky130_fd_sc_hd__clkbuf_1
X_13905_ CPU.registerFile\[31\]\[30\] _07556_ _07557_ CPU.registerFile\[27\]\[30\]
+ _07345_ VGND VGND VPWR VPWR _08318_ sky130_fd_sc_hd__o221a_1
X_17673_ net862 _01961_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16624_ _03987_ VGND VGND VPWR VPWR _02549_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13836_ CPU.registerFile\[21\]\[28\] _07281_ _07521_ CPU.registerFile\[17\]\[28\]
+ _07285_ VGND VGND VPWR VPWR _08251_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_141_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16555_ clknet_1_0__leaf__07219_ VGND VGND VPWR VPWR _03967_ sky130_fd_sc_hd__buf_1
X_10979_ _06191_ VGND VGND VPWR VPWR _02019_ sky130_fd_sc_hd__clkbuf_1
X_13767_ CPU.registerFile\[19\]\[26\] _07383_ _08183_ VGND VGND VPWR VPWR _08184_
+ sky130_fd_sc_hd__o21ai_1
X_15506_ CPU.registerFile\[11\]\[4\] _02861_ VGND VGND VPWR VPWR _03001_ sky130_fd_sc_hd__or2_1
X_12718_ _07198_ _07199_ VGND VGND VPWR VPWR _07200_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16486_ CPU.registerFile\[27\]\[31\] _02928_ _02923_ VGND VGND VPWR VPWR _03954_
+ sky130_fd_sc_hd__o21a_1
X_13698_ CPU.registerFile\[5\]\[24\] _07577_ _08116_ _07638_ VGND VGND VPWR VPWR _08117_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_73_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18225_ net66 _02505_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_15437_ _05029_ VGND VGND VPWR VPWR _02934_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12649_ net1495 _07148_ VGND VGND VPWR VPWR _07151_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14692__797 clknet_1_1__leaf__02684_ VGND VGND VPWR VPWR net829 sky130_fd_sc_hd__inv_2
X_18156_ clknet_leaf_27_clk _02436_ VGND VGND VPWR VPWR CPU.aluIn1\[22\] sky130_fd_sc_hd__dfxtp_4
X_15368_ _02848_ _02857_ _02865_ _08407_ VGND VGND VPWR VPWR _02866_ sky130_fd_sc_hd__o211a_1
X_14391__525 clknet_1_1__leaf__02655_ VGND VGND VPWR VPWR net557 sky130_fd_sc_hd__inv_2
X_17107_ clknet_leaf_23_clk _00040_ VGND VGND VPWR VPWR CPU.cycles\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold305 per_uart.uart0.tx_count16\[2\] VGND VGND VPWR VPWR net1546 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold316 CPU.registerFile\[8\]\[31\] VGND VGND VPWR VPWR net1557 sky130_fd_sc_hd__dlygate4sd3_1
X_18087_ net150 _02367_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15299_ _05405_ VGND VGND VPWR VPWR _02798_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold327 CPU.PC\[22\] VGND VGND VPWR VPWR net1568 sky130_fd_sc_hd__dlygate4sd3_1
X_15044__1111 clknet_1_1__leaf__02721_ VGND VGND VPWR VPWR net1143 sky130_fd_sc_hd__inv_2
Xhold338 CPU.registerFile\[5\]\[9\] VGND VGND VPWR VPWR net1579 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold349 CPU.PC\[7\] VGND VGND VPWR VPWR net1590 sky130_fd_sc_hd__dlygate4sd3_1
X_17038_ net296 _01360_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09860_ _05507_ net1953 _05491_ VGND VGND VPWR VPWR _05508_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__02658_ _02658_ VGND VGND VPWR VPWR clknet_0__02658_ sky130_fd_sc_hd__clkbuf_16
X_08811_ CPU.aluIn1\[2\] _04529_ VGND VGND VPWR VPWR _04531_ sky130_fd_sc_hd__or2_1
X_09791_ _05466_ VGND VGND VPWR VPWR _02529_ sky130_fd_sc_hd__clkbuf_1
Xhold1005 CPU.registerFile\[21\]\[22\] VGND VGND VPWR VPWR net2246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1016 CPU.registerFile\[17\]\[13\] VGND VGND VPWR VPWR net2257 sky130_fd_sc_hd__dlygate4sd3_1
X_08742_ _04459_ _04457_ _04461_ VGND VGND VPWR VPWR _04462_ sky130_fd_sc_hd__o21a_1
Xhold1027 mapped_spi_flash.rcv_data\[0\] VGND VGND VPWR VPWR net2268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1038 CPU.registerFile\[19\]\[6\] VGND VGND VPWR VPWR net2279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 CPU.registerFile\[6\]\[8\] VGND VGND VPWR VPWR net2290 sky130_fd_sc_hd__dlygate4sd3_1
X_08673_ CPU.aluIn1\[14\] VGND VGND VPWR VPWR _04393_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_222 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09225_ _04935_ VGND VGND VPWR VPWR _04936_ sky130_fd_sc_hd__buf_4
XFILLER_0_146_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09156_ _04499_ CPU.Iimm\[3\] _04663_ _04830_ VGND VGND VPWR VPWR _04868_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_79_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09087_ _04799_ VGND VGND VPWR VPWR _02574_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold850 CPU.registerFile\[10\]\[22\] VGND VGND VPWR VPWR net2091 sky130_fd_sc_hd__dlygate4sd3_1
Xhold861 CPU.registerFile\[25\]\[0\] VGND VGND VPWR VPWR net2102 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold872 CPU.registerFile\[25\]\[25\] VGND VGND VPWR VPWR net2113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 CPU.registerFile\[13\]\[18\] VGND VGND VPWR VPWR net2124 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold894 CPU.registerFile\[26\]\[21\] VGND VGND VPWR VPWR net2135 sky130_fd_sc_hd__dlygate4sd3_1
X_10000_ _05555_ net1647 _05558_ VGND VGND VPWR VPWR _05593_ sky130_fd_sc_hd__mux2_1
X_14368__505 clknet_1_1__leaf__02652_ VGND VGND VPWR VPWR net537 sky130_fd_sc_hd__inv_2
X_09989_ _05587_ VGND VGND VPWR VPWR _02452_ sky130_fd_sc_hd__clkbuf_1
X_16638__83 clknet_1_1__leaf__03988_ VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__inv_2
X_11951_ _06742_ VGND VGND VPWR VPWR _01595_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16653__97 clknet_1_1__leaf__03989_ VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__inv_2
X_10902_ _06150_ VGND VGND VPWR VPWR _02055_ sky130_fd_sc_hd__clkbuf_1
X_11882_ net2499 _05729_ _06697_ VGND VGND VPWR VPWR _06706_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__02716_ clknet_0__02716_ VGND VGND VPWR VPWR clknet_1_0__leaf__02716_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_123_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13621_ CPU.registerFile\[6\]\[21\] CPU.registerFile\[7\]\[21\] _07311_ VGND VGND
+ VPWR VPWR _08043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10833_ _06113_ VGND VGND VPWR VPWR _02087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16340_ CPU.registerFile\[18\]\[27\] _02763_ _02770_ _03811_ VGND VGND VPWR VPWR
+ _03812_ sky130_fd_sc_hd__o211a_1
X_13552_ _07411_ _07972_ _07975_ VGND VGND VPWR VPWR _07976_ sky130_fd_sc_hd__or3_1
XFILLER_0_82_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10764_ _05503_ net1605 _06070_ VGND VGND VPWR VPWR _06077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12503_ net2209 _05715_ _07071_ VGND VGND VPWR VPWR _07073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16271_ _02758_ _03742_ _03744_ _05093_ VGND VGND VPWR VPWR _03745_ sky130_fd_sc_hd__a211o_1
X_13483_ _07330_ _07908_ VGND VGND VPWR VPWR _07909_ sky130_fd_sc_hd__or2_1
X_10695_ _06040_ VGND VGND VPWR VPWR _02152_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18010_ net1183 _02290_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_12434_ _07036_ VGND VGND VPWR VPWR _01371_ sky130_fd_sc_hd__clkbuf_1
X_12365_ _05188_ CPU.registerFile\[29\]\[11\] _06999_ VGND VGND VPWR VPWR _07000_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14104_ _08380_ VGND VGND VPWR VPWR _01461_ sky130_fd_sc_hd__clkbuf_1
X_11316_ _05509_ net2318 _06360_ VGND VGND VPWR VPWR _06370_ sky130_fd_sc_hd__mux2_1
X_15084_ _02726_ _02728_ _07181_ VGND VGND VPWR VPWR _02729_ sky130_fd_sc_hd__or3b_1
X_12296_ _06957_ VGND VGND VPWR VPWR _01430_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11247_ _06333_ VGND VGND VPWR VPWR _01893_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11178_ _05507_ net2178 _06288_ VGND VGND VPWR VPWR _06297_ sky130_fd_sc_hd__mux2_1
X_10129_ _05662_ VGND VGND VPWR VPWR _02355_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_143_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15986_ CPU.registerFile\[2\]\[17\] _03227_ _03228_ CPU.registerFile\[3\]\[17\] _03467_
+ VGND VGND VPWR VPWR _03468_ sky130_fd_sc_hd__a221o_1
X_17725_ net914 _02009_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17656_ net845 _01944_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_46_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16607_ _07195_ _03974_ _03975_ _03977_ VGND VGND VPWR VPWR _03978_ sky130_fd_sc_hd__or4_1
X_13819_ net1531 _08018_ _08234_ _08017_ VGND VGND VPWR VPWR _01322_ sky130_fd_sc_hd__o211a_1
X_17587_ net776 _01875_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_840 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_158_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_158_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16469_ _03022_ _03934_ _03935_ _03936_ _03028_ VGND VGND VPWR VPWR _03937_ sky130_fd_sc_hd__o221a_1
X_09010_ _04374_ _04724_ _04726_ VGND VGND VPWR VPWR _04727_ sky130_fd_sc_hd__a21o_1
X_18208_ net49 _02488_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18139_ clknet_leaf_21_clk _02419_ VGND VGND VPWR VPWR CPU.aluIn1\[5\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_14_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16580__52 clknet_1_0__leaf__03969_ VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__inv_2
X_15011__1084 clknet_1_0__leaf__02716_ VGND VGND VPWR VPWR net1116 sky130_fd_sc_hd__inv_2
Xhold102 mapped_spi_flash.cmd_addr\[19\] VGND VGND VPWR VPWR net1343 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 mapped_spi_flash.cmd_addr\[5\] VGND VGND VPWR VPWR net1354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 mapped_spi_flash.cmd_addr\[16\] VGND VGND VPWR VPWR net1365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 mapped_spi_ram.cmd_addr\[4\] VGND VGND VPWR VPWR net1376 sky130_fd_sc_hd__dlygate4sd3_1
X_14317__459 clknet_1_1__leaf__08464_ VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__inv_2
Xhold146 mapped_spi_ram.cmd_addr\[1\] VGND VGND VPWR VPWR net1387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 CPU.mem_wbusy VGND VGND VPWR VPWR net1398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 mapped_spi_ram.cmd_addr\[22\] VGND VGND VPWR VPWR net1409 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09912_ _05305_ VGND VGND VPWR VPWR _05543_ sky130_fd_sc_hd__clkbuf_8
Xhold179 _07137_ VGND VGND VPWR VPWR net1420 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_475 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09843_ _05496_ VGND VGND VPWR VPWR _02507_ sky130_fd_sc_hd__clkbuf_1
X_09774_ _05457_ VGND VGND VPWR VPWR _02537_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08725_ _04444_ VGND VGND VPWR VPWR _04445_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_1_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ _04371_ _04375_ VGND VGND VPWR VPWR _04376_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_1_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_105_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ _04304_ _04289_ _04305_ _04306_ VGND VGND VPWR VPWR _04307_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_37_805 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14675__781 clknet_1_1__leaf__02683_ VGND VGND VPWR VPWR net813 sky130_fd_sc_hd__inv_2
XFILLER_0_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09208_ CPU.PC\[8\] _04919_ VGND VGND VPWR VPWR _04920_ sky130_fd_sc_hd__and2_1
X_10480_ net1400 _05887_ _05851_ _05890_ VGND VGND VPWR VPWR _05891_ sky130_fd_sc_hd__a211o_1
XFILLER_0_134_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09139_ CPU.Jimm\[12\] _04829_ _04831_ VGND VGND VPWR VPWR _04851_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12150_ _05333_ net1906 _06841_ VGND VGND VPWR VPWR _06848_ sky130_fd_sc_hd__mux2_1
X_11101_ _06256_ VGND VGND VPWR VPWR _01962_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12081_ _06811_ VGND VGND VPWR VPWR _01533_ sky130_fd_sc_hd__clkbuf_1
Xhold680 CPU.registerFile\[17\]\[6\] VGND VGND VPWR VPWR net1921 sky130_fd_sc_hd__dlygate4sd3_1
X_14073__347 clknet_1_0__leaf__08367_ VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__inv_2
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold691 CPU.registerFile\[12\]\[30\] VGND VGND VPWR VPWR net1932 sky130_fd_sc_hd__dlygate4sd3_1
X_11032_ _06219_ VGND VGND VPWR VPWR _01994_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_9_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15840_ CPU.registerFile\[22\]\[12\] CPU.registerFile\[23\]\[12\] _02828_ VGND VGND
+ VPWR VPWR _03327_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_125_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15771_ CPU.registerFile\[26\]\[10\] _02861_ VGND VGND VPWR VPWR _03260_ sky130_fd_sc_hd__or2_1
X_12983_ _07308_ VGND VGND VPWR VPWR _07424_ sky130_fd_sc_hd__clkbuf_4
X_17510_ net699 _01798_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_11934_ net2489 _05712_ _06733_ VGND VGND VPWR VPWR _06734_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15043__1110 clknet_1_1__leaf__02721_ VGND VGND VPWR VPWR net1142 sky130_fd_sc_hd__inv_2
X_17441_ net630 _01729_ VGND VGND VPWR VPWR mapped_spi_ram.snd_bitcount\[2\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_2_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_11865_ _06674_ VGND VGND VPWR VPWR _06697_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_28_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14758__856 clknet_1_0__leaf__02691_ VGND VGND VPWR VPWR net888 sky130_fd_sc_hd__inv_2
X_13604_ CPU.registerFile\[28\]\[21\] CPU.registerFile\[24\]\[21\] _04936_ VGND VGND
+ VPWR VPWR _08026_ sky130_fd_sc_hd__mux2_1
X_17372_ net561 _01660_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_10816_ _05555_ net1722 _06069_ VGND VGND VPWR VPWR _06104_ sky130_fd_sc_hd__mux2_1
X_11796_ _06660_ VGND VGND VPWR VPWR _01668_ sky130_fd_sc_hd__clkbuf_1
X_14584_ clknet_1_0__leaf__02664_ VGND VGND VPWR VPWR _02674_ sky130_fd_sc_hd__buf_1
X_16518__186 clknet_1_0__leaf__03963_ VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__inv_2
XFILLER_0_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16323_ CPU.aluIn1\[26\] _07228_ _03778_ _03795_ _06482_ VGND VGND VPWR VPWR _02440_
+ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_41_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13535_ CPU.registerFile\[21\]\[19\] _07502_ _07503_ CPU.registerFile\[17\]\[19\]
+ _07958_ VGND VGND VPWR VPWR _07959_ sky130_fd_sc_hd__o221a_1
XFILLER_0_137_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10747_ _06067_ VGND VGND VPWR VPWR _02127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16254_ _02936_ _03721_ _03728_ _02843_ VGND VGND VPWR VPWR _03729_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13466_ _07306_ _07885_ _07892_ _07703_ VGND VGND VPWR VPWR _07893_ sky130_fd_sc_hd__a31o_1
X_10678_ _04589_ VGND VGND VPWR VPWR _06030_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12417_ _07027_ VGND VGND VPWR VPWR _01379_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_136_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16185_ CPU.registerFile\[1\]\[22\] _02939_ _03661_ _02894_ VGND VGND VPWR VPWR _03662_
+ sky130_fd_sc_hd__a22o_1
X_13397_ CPU.registerFile\[28\]\[14\] CPU.registerFile\[24\]\[14\] _07292_ VGND VGND
+ VPWR VPWR _07826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12348_ _05027_ net2030 _06988_ VGND VGND VPWR VPWR _06991_ sky130_fd_sc_hd__mux2_1
X_12279_ CPU.aluReg\[10\] _06944_ _06924_ VGND VGND VPWR VPWR _06945_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15969_ CPU.registerFile\[5\]\[16\] CPU.registerFile\[4\]\[16\] _03146_ VGND VGND
+ VPWR VPWR _03452_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08510_ CPU.aluIn1\[27\] _04229_ VGND VGND VPWR VPWR _04230_ sky130_fd_sc_hd__and2_1
X_17708_ net897 _01996_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_09490_ net2299 _05188_ _05189_ VGND VGND VPWR VPWR _05190_ sky130_fd_sc_hd__mux2_1
X_17639_ net828 _01927_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_16632__78 clknet_1_0__leaf__03971_ VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__inv_2
XFILLER_0_105_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_156_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15224__134 clknet_1_0__leaf__02753_ VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__inv_2
XFILLER_0_112_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09826_ _05484_ VGND VGND VPWR VPWR _02512_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_107_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09757_ CPU.cycles\[0\] _04687_ _05286_ _05445_ VGND VGND VPWR VPWR _05446_ sky130_fd_sc_hd__a22o_1
X_08708_ _04317_ _04269_ VGND VGND VPWR VPWR _04428_ sky130_fd_sc_hd__nand2b_1
X_09688_ _05365_ _05374_ _05379_ VGND VGND VPWR VPWR _05380_ sky130_fd_sc_hd__or3b_4
XTAP_TAPCELL_ROW_87_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _04230_ _04358_ VGND VGND VPWR VPWR _04359_ sky130_fd_sc_hd__nor2_2
XFILLER_0_96_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11650_ _06573_ VGND VGND VPWR VPWR _06574_ sky130_fd_sc_hd__buf_1
XFILLER_0_37_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10601_ _05967_ VGND VGND VPWR VPWR _05983_ sky130_fd_sc_hd__buf_2
X_11581_ net1378 _06517_ _06509_ _06525_ VGND VGND VPWR VPWR _06526_ sky130_fd_sc_hd__a211o_1
XFILLER_0_107_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13320_ _07254_ _07746_ _07750_ _07268_ VGND VGND VPWR VPWR _07751_ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10532_ _05886_ _04631_ VGND VGND VPWR VPWR _05934_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10463_ CPU.PC\[14\] _04598_ VGND VGND VPWR VPWR _05876_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_118_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13251_ CPU.registerFile\[16\]\[10\] CPU.registerFile\[20\]\[10\] _07258_ VGND VGND
+ VPWR VPWR _07684_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12202_ _06885_ VGND VGND VPWR VPWR _01452_ sky130_fd_sc_hd__clkbuf_1
X_13182_ _07609_ _07616_ _07395_ VGND VGND VPWR VPWR _07617_ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10394_ _05817_ _05823_ VGND VGND VPWR VPWR _05824_ sky130_fd_sc_hd__and2_1
X_12133_ _05150_ net2252 _06830_ VGND VGND VPWR VPWR _06839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15199__111 clknet_1_1__leaf__02751_ VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__inv_2
X_17990_ clknet_leaf_8_clk _02274_ VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16941_ net236 _01267_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_12064_ _06802_ VGND VGND VPWR VPWR _01541_ sky130_fd_sc_hd__clkbuf_1
X_11015_ net2420 _05729_ _06201_ VGND VGND VPWR VPWR _06210_ sky130_fd_sc_hd__mux2_1
X_16872_ _03972_ _04153_ VGND VGND VPWR VPWR _04158_ sky130_fd_sc_hd__nand2_1
X_15823_ CPU.registerFile\[24\]\[12\] _03130_ _02790_ _03309_ VGND VGND VPWR VPWR
+ _03310_ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15754_ CPU.registerFile\[14\]\[10\] _02889_ VGND VGND VPWR VPWR _03243_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12966_ CPU.registerFile\[29\]\[2\] _07403_ _07404_ CPU.registerFile\[25\]\[2\] _07250_
+ VGND VGND VPWR VPWR _07407_ sky130_fd_sc_hd__o221a_1
X_15010__1083 clknet_1_0__leaf__02716_ VGND VGND VPWR VPWR net1115 sky130_fd_sc_hd__inv_2
X_11917_ CPU.registerFile\[11\]\[19\] _05696_ _06722_ VGND VGND VPWR VPWR _06725_
+ sky130_fd_sc_hd__mux2_1
X_14346__485 clknet_1_1__leaf__08467_ VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__inv_2
X_15685_ _03171_ _03175_ _03138_ VGND VGND VPWR VPWR _03176_ sky130_fd_sc_hd__a21o_1
XANTENNA_350 _05380_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12897_ _05283_ VGND VGND VPWR VPWR _07339_ sky130_fd_sc_hd__buf_6
XANTENNA_361 _07356_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_372 _07233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17424_ net613 net1425 VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_383 _05272_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11848_ _06688_ VGND VGND VPWR VPWR _01644_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_394 _07621_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13984__267 clknet_1_0__leaf__08358_ VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__inv_2
XFILLER_0_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ net544 _01643_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11779_ _05008_ net1994 _06650_ VGND VGND VPWR VPWR _06652_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16306_ CPU.registerFile\[28\]\[26\] CPU.registerFile\[24\]\[26\] _02881_ VGND VGND
+ VPWR VPWR _03779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13518_ CPU.registerFile\[13\]\[18\] _07482_ _07420_ CPU.registerFile\[9\]\[18\]
+ _07249_ VGND VGND VPWR VPWR _07943_ sky130_fd_sc_hd__o221a_1
X_17286_ net475 _01574_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload11 clknet_leaf_14_clk VGND VGND VPWR VPWR clkload11/Y sky130_fd_sc_hd__clkinv_4
X_16237_ CPU.registerFile\[29\]\[24\] _02918_ VGND VGND VPWR VPWR _03712_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_151_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13449_ _07570_ _07875_ VGND VGND VPWR VPWR _07876_ sky130_fd_sc_hd__or2_1
Xclkload22 clknet_leaf_3_clk VGND VGND VPWR VPWR clkload22/Y sky130_fd_sc_hd__inv_6
Xclkload33 clknet_1_0__leaf__02753_ VGND VGND VPWR VPWR clkload33/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload44 clknet_1_0__leaf__02723_ VGND VGND VPWR VPWR clkload44/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload55 clknet_1_0__leaf__02701_ VGND VGND VPWR VPWR clkload55/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16168_ CPU.registerFile\[27\]\[22\] CPU.registerFile\[31\]\[22\] _02852_ VGND VGND
+ VPWR VPWR _03645_ sky130_fd_sc_hd__mux2_1
Xclkload66 clknet_1_1__leaf__02685_ VGND VGND VPWR VPWR clkload66/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload77 clknet_1_1__leaf__02667_ VGND VGND VPWR VPWR clkload77/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload88 clknet_1_1__leaf__02656_ VGND VGND VPWR VPWR clkload88/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload99 clknet_1_1__leaf__08430_ VGND VGND VPWR VPWR clkload99/Y sky130_fd_sc_hd__clkinvlp_4
X_15119_ clknet_1_1__leaf__02720_ VGND VGND VPWR VPWR _02743_ sky130_fd_sc_hd__buf_1
XFILLER_0_2_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14056__331 clknet_1_0__leaf__08366_ VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_54_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08990_ _04491_ VGND VGND VPWR VPWR _04708_ sky130_fd_sc_hd__clkbuf_4
X_16099_ _02949_ _03574_ _03577_ VGND VGND VPWR VPWR _03578_ sky130_fd_sc_hd__or3_2
X_14511__633 clknet_1_1__leaf__02667_ VGND VGND VPWR VPWR net665 sky130_fd_sc_hd__inv_2
XFILLER_0_11_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09611_ _05305_ VGND VGND VPWR VPWR _05306_ sky130_fd_sc_hd__clkbuf_8
X_09542_ _04885_ _05238_ VGND VGND VPWR VPWR _05239_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_92_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09473_ _04744_ _05172_ _04636_ VGND VGND VPWR VPWR _05173_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_102_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload5 clknet_leaf_26_clk VGND VGND VPWR VPWR clkload5/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_144_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14787__882 clknet_1_0__leaf__02694_ VGND VGND VPWR VPWR net914 sky130_fd_sc_hd__inv_2
XFILLER_0_112_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14486__610 clknet_1_1__leaf__02665_ VGND VGND VPWR VPWR net642 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_89_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09809_ net1705 _05209_ _05474_ VGND VGND VPWR VPWR _05476_ sky130_fd_sc_hd__mux2_1
X_12820_ _05336_ VGND VGND VPWR VPWR _07263_ sky130_fd_sc_hd__buf_4
XFILLER_0_97_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14226__401 clknet_1_0__leaf__08432_ VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__inv_2
XFILLER_0_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11702_ mapped_spi_ram.rcv_data\[10\] _06601_ VGND VGND VPWR VPWR _06605_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15470_ _02914_ _02964_ _02965_ VGND VGND VPWR VPWR _02966_ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12682_ _07168_ net1429 VGND VGND VPWR VPWR _00033_ sky130_fd_sc_hd__nor2_1
X_11633_ _06550_ _06560_ VGND VGND VPWR VPWR _06561_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17140_ net364 _01428_ VGND VGND VPWR VPWR CPU.aluReg\[4\] sky130_fd_sc_hd__dfxtp_1
X_11564_ _06512_ _05889_ VGND VGND VPWR VPWR _06513_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13303_ _07411_ _07731_ _07734_ VGND VGND VPWR VPWR _07735_ sky130_fd_sc_hd__or3_1
X_17071_ net329 _01393_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_10515_ net1384 _05887_ _05856_ _05920_ VGND VGND VPWR VPWR _05921_ sky130_fd_sc_hd__a211o_1
X_14283_ _08456_ _08458_ _08460_ _08461_ _06482_ VGND VGND VPWR VPWR _01559_ sky130_fd_sc_hd__o311a_1
X_11495_ _05551_ net2472 _06455_ VGND VGND VPWR VPWR _06465_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_133_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16022_ CPU.registerFile\[13\]\[18\] _03123_ VGND VGND VPWR VPWR _03503_ sky130_fd_sc_hd__or2_1
X_13234_ _07398_ _07666_ _07667_ VGND VGND VPWR VPWR _07668_ sky130_fd_sc_hd__o21a_1
X_10446_ net1401 _05849_ _05862_ _05855_ VGND VGND VPWR VPWR _02222_ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__02660_ clknet_0__02660_ VGND VGND VPWR VPWR clknet_1_1__leaf__02660_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_110_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__02691_ _02691_ VGND VGND VPWR VPWR clknet_0__02691_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_21_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13165_ _07397_ _07593_ _07600_ _07424_ VGND VGND VPWR VPWR _07601_ sky130_fd_sc_hd__a31o_2
X_10377_ _05810_ VGND VGND VPWR VPWR _02240_ sky130_fd_sc_hd__clkbuf_1
X_12116_ _06818_ VGND VGND VPWR VPWR _06830_ sky130_fd_sc_hd__buf_4
X_17973_ net1161 _02257_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_13096_ CPU.registerFile\[18\]\[6\] CPU.registerFile\[22\]\[6\] _07240_ VGND VGND
+ VPWR VPWR _07533_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12047_ _06793_ VGND VGND VPWR VPWR _01549_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_148_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16855_ net1797 per_uart.rx_data\[6\] _04139_ VGND VGND VPWR VPWR _04146_ sky130_fd_sc_hd__mux2_1
X_15806_ CPU.registerFile\[18\]\[11\] _02832_ _02835_ CPU.registerFile\[19\]\[11\]
+ _03074_ VGND VGND VPWR VPWR _03294_ sky130_fd_sc_hd__o221a_1
XFILLER_0_88_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16786_ _04052_ _04978_ _08453_ VGND VGND VPWR VPWR _04098_ sky130_fd_sc_hd__or3b_1
X_13998_ clknet_1_0__leaf__07223_ VGND VGND VPWR VPWR _08360_ sky130_fd_sc_hd__buf_1
X_15737_ CPU.registerFile\[1\]\[10\] _03030_ _03225_ _03028_ VGND VGND VPWR VPWR _03226_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15253__160 clknet_1_1__leaf__02756_ VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__inv_2
X_12949_ CPU.registerFile\[5\]\[2\] _04987_ _07389_ _07368_ VGND VGND VPWR VPWR _07390_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_888 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15668_ CPU.registerFile\[14\]\[8\] CPU.registerFile\[10\]\[8\] _03082_ VGND VGND
+ VPWR VPWR _03159_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_180 _07555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_191 _07841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17407_ net596 _01695_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15599_ CPU.registerFile\[30\]\[6\] CPU.registerFile\[26\]\[6\] _02787_ VGND VGND
+ VPWR VPWR _03092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17338_ net527 _01626_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload100 clknet_1_0__leaf__08429_ VGND VGND VPWR VPWR clkload100/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_114_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18370__29 VGND VGND VPWR VPWR _18370__29/HI net29 sky130_fd_sc_hd__conb_1
Xclkload111 clknet_1_0__leaf__07219_ VGND VGND VPWR VPWR clkload111/X sky130_fd_sc_hd__clkbuf_8
X_17269_ net459 _01557_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__08434_ clknet_0__08434_ VGND VGND VPWR VPWR clknet_1_1__leaf__08434_
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_0__08465_ _08465_ VGND VGND VPWR VPWR clknet_0__08465_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__08365_ clknet_0__08365_ VGND VGND VPWR VPWR clknet_1_1__leaf__08365_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08973_ mapped_spi_ram.rcv_data\[6\] _04689_ _04691_ mapped_spi_flash.rcv_data\[6\]
+ VGND VGND VPWR VPWR _04692_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__02680_ clknet_0__02680_ VGND VGND VPWR VPWR clknet_1_0__leaf__02680_
+ sky130_fd_sc_hd__clkbuf_16
X_09525_ _05220_ _05222_ _04708_ VGND VGND VPWR VPWR _05223_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_84_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13967__251 clknet_1_0__leaf__08357_ VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__inv_2
X_09456_ _04325_ _04698_ _04210_ _04262_ VGND VGND VPWR VPWR _05157_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09387_ _05091_ VGND VGND VPWR VPWR _02566_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14221__397 clknet_1_0__leaf__08431_ VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_115_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10300_ _05769_ VGND VGND VPWR VPWR _02291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11280_ CPU.registerFile\[9\]\[7\] _05721_ _06346_ VGND VGND VPWR VPWR _06351_ sky130_fd_sc_hd__mux2_1
X_10231_ _05730_ VGND VGND VPWR VPWR _02321_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10162_ net2032 _05683_ _05671_ VGND VGND VPWR VPWR _05684_ sky130_fd_sc_hd__mux2_1
X_14989__1064 clknet_1_0__leaf__02714_ VGND VGND VPWR VPWR net1096 sky130_fd_sc_hd__inv_2
X_10093_ _05643_ VGND VGND VPWR VPWR _02372_ sky130_fd_sc_hd__clkbuf_1
X_13921_ CPU.registerFile\[19\]\[31\] _07618_ _08332_ _07417_ _07278_ VGND VGND VPWR
+ VPWR _08333_ sky130_fd_sc_hd__o221a_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13852_ CPU.registerFile\[6\]\[29\] CPU.registerFile\[7\]\[29\] _07641_ VGND VGND
+ VPWR VPWR _08266_ sky130_fd_sc_hd__mux2_1
X_12803_ CPU.registerFile\[16\]\[0\] CPU.registerFile\[20\]\[0\] _07240_ VGND VGND
+ VPWR VPWR _07246_ sky130_fd_sc_hd__mux2_1
X_13783_ CPU.registerFile\[14\]\[26\] CPU.registerFile\[10\]\[26\] _07476_ VGND VGND
+ VPWR VPWR _08200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10995_ _06199_ VGND VGND VPWR VPWR _02011_ sky130_fd_sc_hd__clkbuf_1
X_18310_ clknet_leaf_16_clk _02590_ VGND VGND VPWR VPWR CPU.PC\[10\] sky130_fd_sc_hd__dfxtp_1
X_15522_ CPU.registerFile\[25\]\[4\] CPU.registerFile\[29\]\[4\] _02851_ VGND VGND
+ VPWR VPWR _03017_ sky130_fd_sc_hd__mux2_1
X_12734_ _07212_ VGND VGND VPWR VPWR _01259_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18241_ net82 _02521_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_15453_ CPU.registerFile\[20\]\[2\] CPU.registerFile\[21\]\[2\] _08395_ VGND VGND
+ VPWR VPWR _02950_ sky130_fd_sc_hd__mux2_1
X_12665_ net1485 _07158_ VGND VGND VPWR VPWR _00025_ sky130_fd_sc_hd__xor2_1
XFILLER_0_26_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18172_ net203 _02452_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11616_ _06469_ _06471_ _06486_ net1930 VGND VGND VPWR VPWR _06547_ sky130_fd_sc_hd__o31a_1
XFILLER_0_154_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15384_ CPU.registerFile\[28\]\[1\] CPU.registerFile\[24\]\[1\] _02881_ VGND VGND
+ VPWR VPWR _02882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12596_ _04292_ _05134_ _04653_ VGND VGND VPWR VPWR _07122_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_154_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17123_ clknet_leaf_17_clk _00025_ VGND VGND VPWR VPWR CPU.cycles\[19\] sky130_fd_sc_hd__dfxtp_1
X_14458__586 clknet_1_1__leaf__02661_ VGND VGND VPWR VPWR net618 sky130_fd_sc_hd__inv_2
X_11547_ net1345 _06495_ _06500_ _06006_ VGND VGND VPWR VPWR _01756_ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17054_ net312 _01376_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[16\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__02712_ clknet_0__02712_ VGND VGND VPWR VPWR clknet_1_1__leaf__02712_
+ sky130_fd_sc_hd__clkbuf_16
Xhold509 per_uart.d_in_uart\[2\] VGND VGND VPWR VPWR net1750 sky130_fd_sc_hd__dlygate4sd3_1
X_14266_ _04724_ _04765_ _04788_ _08444_ VGND VGND VPWR VPWR _08445_ sky130_fd_sc_hd__or4_1
XFILLER_0_40_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14196__374 clknet_1_1__leaf__08429_ VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__inv_2
X_11478_ _06456_ VGND VGND VPWR VPWR _01785_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16005_ _03482_ _03486_ _03252_ VGND VGND VPWR VPWR _03487_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13217_ CPU.registerFile\[23\]\[9\] _07382_ _07649_ _07650_ _07288_ VGND VGND VPWR
+ VPWR _07651_ sky130_fd_sc_hd__o221a_1
Xclkbuf_0__02743_ _02743_ VGND VGND VPWR VPWR clknet_0__02743_ sky130_fd_sc_hd__clkbuf_16
X_10429_ _05842_ VGND VGND VPWR VPWR _05849_ sky130_fd_sc_hd__buf_2
XFILLER_0_110_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13148_ _07302_ VGND VGND VPWR VPWR _07584_ sky130_fd_sc_hd__buf_8
Xclkbuf_0__02674_ _02674_ VGND VGND VPWR VPWR clknet_0__02674_ sky130_fd_sc_hd__clkbuf_16
X_13079_ CPU.registerFile\[15\]\[5\] _07276_ _07277_ CPU.registerFile\[11\]\[5\] _07278_
+ VGND VGND VPWR VPWR _07517_ sky130_fd_sc_hd__o221a_1
X_17956_ net1144 _02240_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[1\] sky130_fd_sc_hd__dfxtp_1
Xhold1209 CPU.registerFile\[1\]\[20\] VGND VGND VPWR VPWR net2450 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_29_Left_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_146_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16907_ _04631_ _04635_ _04181_ _06468_ VGND VGND VPWR VPWR _04182_ sky130_fd_sc_hd__and4b_2
X_17887_ net1076 _02171_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14623__734 clknet_1_0__leaf__02678_ VGND VGND VPWR VPWR net766 sky130_fd_sc_hd__inv_2
X_16838_ _05816_ _04135_ VGND VGND VPWR VPWR _04136_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16769_ _03995_ _05035_ _07132_ VGND VGND VPWR VPWR _04084_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_66_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09310_ _04448_ _04806_ VGND VGND VPWR VPWR _05018_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09241_ _04908_ _04951_ VGND VGND VPWR VPWR _04952_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_1_Left_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_38_Left_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09172_ CPU.PC\[7\] CPU.Bimm\[7\] _04819_ VGND VGND VPWR VPWR _04884_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08956_ _04367_ _04224_ _04365_ VGND VGND VPWR VPWR _04675_ sky130_fd_sc_hd__or3_1
X_08887_ _04565_ _04566_ _04605_ _04506_ VGND VGND VPWR VPWR _04607_ sky130_fd_sc_hd__a31o_1
XFILLER_0_98_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14899__983 clknet_1_0__leaf__02705_ VGND VGND VPWR VPWR net1015 sky130_fd_sc_hd__inv_2
XFILLER_0_79_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14598__711 clknet_1_1__leaf__02676_ VGND VGND VPWR VPWR net743 sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__02663_ clknet_0__02663_ VGND VGND VPWR VPWR clknet_1_0__leaf__02663_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09508_ _04974_ _05195_ _05197_ _04955_ _05206_ VGND VGND VPWR VPWR _05207_ sky130_fd_sc_hd__o221ai_4
X_10780_ _06085_ VGND VGND VPWR VPWR _02112_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09439_ CPU.aluIn1\[13\] _04259_ _04698_ VGND VGND VPWR VPWR _05141_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12450_ _07044_ VGND VGND VPWR VPWR _01363_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_10_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11401_ _06415_ VGND VGND VPWR VPWR _01821_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12381_ _05381_ net2180 _06999_ VGND VGND VPWR VPWR _07008_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_80 _05208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_91 _05306_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14120_ _05172_ VGND VGND VPWR VPWR _08389_ sky130_fd_sc_hd__inv_2
X_11332_ _06378_ VGND VGND VPWR VPWR _01853_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11263_ CPU.registerFile\[9\]\[15\] _05704_ _06335_ VGND VGND VPWR VPWR _06342_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13002_ CPU.registerFile\[14\]\[3\] CPU.registerFile\[10\]\[3\] _07274_ VGND VGND
+ VPWR VPWR _07442_ sky130_fd_sc_hd__mux2_1
X_10214_ _05252_ VGND VGND VPWR VPWR _05719_ sky130_fd_sc_hd__clkbuf_4
X_11194_ _06305_ VGND VGND VPWR VPWR _01918_ sky130_fd_sc_hd__clkbuf_1
X_10145_ _05672_ VGND VGND VPWR VPWR _02349_ sky130_fd_sc_hd__clkbuf_1
X_17810_ net999 _02094_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17741_ net930 _02025_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[27\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_128_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10076_ net1664 _04696_ _05633_ VGND VGND VPWR VPWR _05635_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13904_ _07351_ _08316_ VGND VGND VPWR VPWR _08317_ sky130_fd_sc_hd__or2_1
X_17672_ net861 _01960_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14884_ clknet_1_1__leaf__02697_ VGND VGND VPWR VPWR _02704_ sky130_fd_sc_hd__buf_1
X_16623_ per_uart.uart0.uart_rxd2 net1825 _03979_ VGND VGND VPWR VPWR _03987_ sky130_fd_sc_hd__mux2_1
X_13835_ CPU.registerFile\[16\]\[28\] CPU.registerFile\[20\]\[28\] _07785_ VGND VGND
+ VPWR VPWR _08250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_27_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_141_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13766_ CPU.registerFile\[23\]\[26\] _07382_ _08182_ _07418_ _07288_ VGND VGND VPWR
+ VPWR _08183_ sky130_fd_sc_hd__o221a_1
X_10978_ net1672 _05691_ _06190_ VGND VGND VPWR VPWR _06191_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__08368_ clknet_0__08368_ VGND VGND VPWR VPWR clknet_1_0__leaf__08368_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15505_ CPU.registerFile\[9\]\[4\] CPU.registerFile\[13\]\[4\] _02999_ VGND VGND
+ VPWR VPWR _03000_ sky130_fd_sc_hd__mux2_1
X_12717_ per_uart.uart0.tx_bitcount\[2\] per_uart.uart0.tx_bitcount\[0\] per_uart.uart0.tx_bitcount\[1\]
+ per_uart.uart0.tx_bitcount\[3\] VGND VGND VPWR VPWR _07199_ sky130_fd_sc_hd__and4bb_1
X_16485_ CPU.registerFile\[31\]\[31\] _03072_ VGND VGND VPWR VPWR _03953_ sky130_fd_sc_hd__or2_1
X_13697_ CPU.registerFile\[4\]\[24\] _07374_ VGND VGND VPWR VPWR _08116_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18224_ net65 _02504_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_61_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15436_ _08411_ _02917_ _02932_ _08408_ VGND VGND VPWR VPWR _02933_ sky130_fd_sc_hd__o211a_1
X_12648_ CPU.cycles\[12\] _07148_ VGND VGND VPWR VPWR _07150_ sky130_fd_sc_hd__and2_1
XFILLER_0_155_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14811__904 clknet_1_0__leaf__02696_ VGND VGND VPWR VPWR net936 sky130_fd_sc_hd__inv_2
X_14204__381 clknet_1_0__leaf__08430_ VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__inv_2
X_18155_ clknet_leaf_22_clk _02435_ VGND VGND VPWR VPWR CPU.aluIn1\[21\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_25_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15367_ _02858_ _02859_ _02863_ _02864_ VGND VGND VPWR VPWR _02865_ sky130_fd_sc_hd__a211o_1
X_12579_ CPU.registerFile\[4\]\[6\] _05305_ _07107_ VGND VGND VPWR VPWR _07113_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17106_ clknet_leaf_23_clk _00037_ VGND VGND VPWR VPWR CPU.cycles\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14318_ clknet_1_0__leaf__08433_ VGND VGND VPWR VPWR _08465_ sky130_fd_sc_hd__buf_1
X_18086_ net149 _02366_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[16\] sky130_fd_sc_hd__dfxtp_1
Xhold306 CPU.registerFile\[5\]\[10\] VGND VGND VPWR VPWR net1547 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15298_ _02796_ VGND VGND VPWR VPWR _02797_ sky130_fd_sc_hd__buf_4
Xhold317 CPU.registerFile\[5\]\[7\] VGND VGND VPWR VPWR net1558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 CPU.PC\[14\] VGND VGND VPWR VPWR net1569 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12751__204 clknet_1_0__leaf__07221_ VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__inv_2
XFILLER_0_1_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17037_ net295 _01359_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[31\] sky130_fd_sc_hd__dfxtp_1
Xhold339 CPU.registerFile\[16\]\[30\] VGND VGND VPWR VPWR net1580 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_471 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08810_ CPU.aluIn1\[2\] _04529_ VGND VGND VPWR VPWR _04530_ sky130_fd_sc_hd__nand2_1
Xclkbuf_0__02657_ _02657_ VGND VGND VPWR VPWR clknet_0__02657_ sky130_fd_sc_hd__clkbuf_16
X_09790_ net1923 _05027_ _05463_ VGND VGND VPWR VPWR _05466_ sky130_fd_sc_hd__mux2_1
Xhold1006 CPU.registerFile\[25\]\[5\] VGND VGND VPWR VPWR net2247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1017 CPU.registerFile\[23\]\[20\] VGND VGND VPWR VPWR net2258 sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ _04460_ _04348_ VGND VGND VPWR VPWR _04461_ sky130_fd_sc_hd__nand2_2
Xhold1028 CPU.registerFile\[13\]\[9\] VGND VGND VPWR VPWR net2269 sky130_fd_sc_hd__dlygate4sd3_1
X_17939_ net1128 _02223_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[19\] sky130_fd_sc_hd__dfxtp_1
Xhold1039 CPU.registerFile\[31\]\[11\] VGND VGND VPWR VPWR net2280 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08672_ _04391_ _04255_ VGND VGND VPWR VPWR _04392_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_814 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_18_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_46_Left_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_908 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_118_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09224_ mapped_spi_ram.rcv_data\[14\] net18 _04618_ mapped_spi_flash.rcv_data\[14\]
+ VGND VGND VPWR VPWR _04935_ sky130_fd_sc_hd__a22oi_4
X_14988__1063 clknet_1_0__leaf__02714_ VGND VGND VPWR VPWR net1095 sky130_fd_sc_hd__inv_2
XFILLER_0_17_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09155_ CPU.PC\[4\] _04866_ VGND VGND VPWR VPWR _04867_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09086_ net2207 _04798_ _04668_ VGND VGND VPWR VPWR _04799_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold840 CPU.registerFile\[24\]\[12\] VGND VGND VPWR VPWR net2081 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_55_Left_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold851 CPU.registerFile\[27\]\[26\] VGND VGND VPWR VPWR net2092 sky130_fd_sc_hd__dlygate4sd3_1
Xhold862 CPU.registerFile\[3\]\[7\] VGND VGND VPWR VPWR net2103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 CPU.registerFile\[7\]\[0\] VGND VGND VPWR VPWR net2114 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold884 CPU.registerFile\[3\]\[4\] VGND VGND VPWR VPWR net2125 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold895 CPU.registerFile\[22\]\[7\] VGND VGND VPWR VPWR net2136 sky130_fd_sc_hd__dlygate4sd3_1
X_09988_ _05543_ net2495 _05581_ VGND VGND VPWR VPWR _05587_ sky130_fd_sc_hd__mux2_1
X_14907__990 clknet_1_1__leaf__02706_ VGND VGND VPWR VPWR net1022 sky130_fd_sc_hd__inv_2
X_08939_ _04658_ VGND VGND VPWR VPWR _04659_ sky130_fd_sc_hd__buf_4
X_15193__106 clknet_1_0__leaf__02750_ VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_150_Right_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11950_ CPU.registerFile\[11\]\[3\] _05729_ _06733_ VGND VGND VPWR VPWR _06742_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10901_ net1649 _05683_ _06143_ VGND VGND VPWR VPWR _06150_ sky130_fd_sc_hd__mux2_1
X_11881_ _06705_ VGND VGND VPWR VPWR _01628_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__02715_ clknet_0__02715_ VGND VGND VPWR VPWR clknet_1_0__leaf__02715_
+ sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_64_Left_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_123_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13620_ CPU.registerFile\[1\]\[21\] _07256_ _08041_ _07368_ VGND VGND VPWR VPWR _08042_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_123_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10832_ net1709 _05683_ _06106_ VGND VGND VPWR VPWR _06113_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13551_ CPU.registerFile\[11\]\[19\] _07363_ _07974_ VGND VGND VPWR VPWR _07975_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_109_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10763_ _06076_ VGND VGND VPWR VPWR _02120_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12502_ _07072_ VGND VGND VPWR VPWR _01339_ sky130_fd_sc_hd__clkbuf_1
X_16270_ CPU.registerFile\[25\]\[25\] _05406_ _02779_ _03743_ VGND VGND VPWR VPWR
+ _03744_ sky130_fd_sc_hd__o211a_1
X_13482_ CPU.registerFile\[18\]\[17\] CPU.registerFile\[22\]\[17\] _07314_ VGND VGND
+ VPWR VPWR _07908_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10694_ _05501_ net1761 _06034_ VGND VGND VPWR VPWR _06040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12433_ _05188_ net2280 _07035_ VGND VGND VPWR VPWR _07036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15152_ clknet_1_0__leaf__02720_ VGND VGND VPWR VPWR _02746_ sky130_fd_sc_hd__buf_1
X_14652__760 clknet_1_0__leaf__02681_ VGND VGND VPWR VPWR net792 sky130_fd_sc_hd__inv_2
X_12364_ _06976_ VGND VGND VPWR VPWR _06999_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_73_Left_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14103_ _08379_ _05363_ _00000_ VGND VGND VPWR VPWR _08380_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11315_ _06369_ VGND VGND VPWR VPWR _01861_ sky130_fd_sc_hd__clkbuf_1
X_15083_ per_uart.uart0.enable16_counter\[2\] _07180_ VGND VGND VPWR VPWR _02728_
+ sky130_fd_sc_hd__and2_1
X_12295_ net2484 _06956_ _06861_ VGND VGND VPWR VPWR _06957_ sky130_fd_sc_hd__mux2_1
X_11246_ CPU.registerFile\[9\]\[23\] _05687_ _06324_ VGND VGND VPWR VPWR _06333_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11177_ _06296_ VGND VGND VPWR VPWR _01926_ sky130_fd_sc_hd__clkbuf_1
X_14050__326 clknet_1_0__leaf__08365_ VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__inv_2
X_10128_ net2063 _05333_ _05655_ VGND VGND VPWR VPWR _05662_ sky130_fd_sc_hd__mux2_1
X_15985_ CPU.registerFile\[7\]\[17\] _02898_ _02887_ _03466_ VGND VGND VPWR VPWR _03467_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_143_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17724_ net913 _02008_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_10059_ net2212 _05333_ _05618_ VGND VGND VPWR VPWR _05625_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_82_Left_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17655_ net844 _01943_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_46_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16606_ net2 _03976_ VGND VGND VPWR VPWR _03977_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_34_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13818_ _07394_ _08219_ _08233_ _08015_ VGND VGND VPWR VPWR _08234_ sky130_fd_sc_hd__a211o_1
XFILLER_0_86_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17586_ net775 _01874_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13749_ CPU.registerFile\[14\]\[25\] CPU.registerFile\[6\]\[25\] _04648_ VGND VGND
+ VPWR VPWR _08167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_158_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_158_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14735__835 clknet_1_0__leaf__02689_ VGND VGND VPWR VPWR net867 sky130_fd_sc_hd__inv_2
X_16468_ CPU.registerFile\[20\]\[31\] _02855_ _03026_ VGND VGND VPWR VPWR _03936_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_362 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15419_ _02914_ _02915_ _02848_ VGND VGND VPWR VPWR _02916_ sky130_fd_sc_hd__a21o_1
X_18207_ net48 _02487_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_16399_ CPU.registerFile\[21\]\[29\] CPU.registerFile\[23\]\[29\] _02769_ VGND VGND
+ VPWR VPWR _03869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_91_Left_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18138_ clknet_leaf_27_clk _02418_ VGND VGND VPWR VPWR CPU.aluIn1\[4\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_14_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold103 mapped_spi_ram.rcv_bitcount\[3\] VGND VGND VPWR VPWR net1344 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold114 CPU.cycles\[5\] VGND VGND VPWR VPWR net1355 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18069_ net132 _02349_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_87 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold125 mapped_spi_flash.cmd_addr\[9\] VGND VGND VPWR VPWR net1366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_7_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_8
Xhold136 mapped_spi_flash.cmd_addr\[13\] VGND VGND VPWR VPWR net1377 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 mapped_spi_ram.cmd_addr\[5\] VGND VGND VPWR VPWR net1388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 mapped_spi_flash.cmd_addr\[15\] VGND VGND VPWR VPWR net1399 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ _05542_ VGND VGND VPWR VPWR _02485_ sky130_fd_sc_hd__clkbuf_1
Xhold169 per_uart.uart0.txd_reg\[7\] VGND VGND VPWR VPWR net1410 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__02709_ _02709_ VGND VGND VPWR VPWR clknet_0__02709_ sky130_fd_sc_hd__clkbuf_16
X_09842_ _05495_ net2347 _05491_ VGND VGND VPWR VPWR _05496_ sky130_fd_sc_hd__mux2_1
X_09773_ net2216 _04748_ _05452_ VGND VGND VPWR VPWR _05457_ sky130_fd_sc_hd__mux2_1
X_14781__877 clknet_1_0__leaf__02693_ VGND VGND VPWR VPWR net909 sky130_fd_sc_hd__inv_2
X_08724_ _04337_ _04250_ VGND VGND VPWR VPWR _04444_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08655_ _04370_ _04222_ _04368_ _04374_ VGND VGND VPWR VPWR _04375_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_1_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08586_ CPU.aluIn1\[2\] net1292 VGND VGND VPWR VPWR _04306_ sky130_fd_sc_hd__nand2_2
XFILLER_0_138_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14027__306 clknet_1_1__leaf__08362_ VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__inv_2
XFILLER_0_138_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09207_ CPU.PC\[7\] CPU.PC\[6\] _04918_ VGND VGND VPWR VPWR _04919_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_20_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09138_ _04848_ _04849_ VGND VGND VPWR VPWR _04850_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09069_ _04504_ VGND VGND VPWR VPWR _04782_ sky130_fd_sc_hd__buf_2
X_11100_ net2500 _05677_ _06252_ VGND VGND VPWR VPWR _06256_ sky130_fd_sc_hd__mux2_1
X_12080_ _05306_ net1794 _06805_ VGND VGND VPWR VPWR _06811_ sky130_fd_sc_hd__mux2_1
Xhold670 CPU.registerFile\[23\]\[16\] VGND VGND VPWR VPWR net1911 sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 CPU.registerFile\[31\]\[5\] VGND VGND VPWR VPWR net1922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 CPU.registerFile\[3\]\[31\] VGND VGND VPWR VPWR net1933 sky130_fd_sc_hd__dlygate4sd3_1
X_11031_ net1878 _05677_ _06215_ VGND VGND VPWR VPWR _06219_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15201__113 clknet_1_1__leaf__02751_ VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_125_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15770_ CPU.registerFile\[28\]\[10\] CPU.registerFile\[24\]\[10\] _02918_ VGND VGND
+ VPWR VPWR _03259_ sky130_fd_sc_hd__mux2_1
X_12982_ _07411_ _07416_ _07422_ VGND VGND VPWR VPWR _07423_ sky130_fd_sc_hd__or3_2
X_11933_ _06710_ VGND VGND VPWR VPWR _06733_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17440_ net629 _01728_ VGND VGND VPWR VPWR mapped_spi_ram.snd_bitcount\[1\] sky130_fd_sc_hd__dfxtp_1
X_11864_ _06696_ VGND VGND VPWR VPWR _01636_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ _08021_ _08024_ _07405_ VGND VGND VPWR VPWR _08025_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17371_ net560 _01659_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_10815_ _06103_ VGND VGND VPWR VPWR _02095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11795_ _05170_ net1986 _06650_ VGND VGND VPWR VPWR _06660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16322_ _08411_ _03786_ _03794_ _07308_ VGND VGND VPWR VPWR _03795_ sky130_fd_sc_hd__a31o_1
X_13534_ _07245_ _07957_ VGND VGND VPWR VPWR _07958_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_41_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10746_ _05553_ net1678 _06033_ VGND VGND VPWR VPWR _06067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16253_ _05010_ _03724_ _03727_ VGND VGND VPWR VPWR _03728_ sky130_fd_sc_hd__or3_2
X_13465_ _07231_ _07888_ _07891_ VGND VGND VPWR VPWR _07892_ sky130_fd_sc_hd__or3_1
XFILLER_0_82_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10677_ _06029_ VGND VGND VPWR VPWR _02159_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12416_ _05027_ net2231 _07024_ VGND VGND VPWR VPWR _07027_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_136_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16184_ CPU.registerFile\[5\]\[22\] CPU.registerFile\[4\]\[22\] _03146_ VGND VGND
+ VPWR VPWR _03661_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_136_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13396_ _07519_ _07823_ _07824_ VGND VGND VPWR VPWR _07825_ sky130_fd_sc_hd__o21a_1
XFILLER_0_51_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12347_ _06990_ VGND VGND VPWR VPWR _01412_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12278_ CPU.aluIn1\[10\] _06943_ _06927_ VGND VGND VPWR VPWR _06944_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11229_ _06323_ VGND VGND VPWR VPWR _06324_ sky130_fd_sc_hd__buf_4
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14987__1062 clknet_1_0__leaf__02714_ VGND VGND VPWR VPWR net1094 sky130_fd_sc_hd__inv_2
X_15968_ CPU.registerFile\[2\]\[16\] _03143_ _02980_ CPU.registerFile\[3\]\[16\] _03144_
+ VGND VGND VPWR VPWR _03451_ sky130_fd_sc_hd__a221o_1
X_17707_ net896 _01995_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_15899_ CPU.registerFile\[7\]\[14\] _03317_ VGND VGND VPWR VPWR _03384_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17638_ net827 _01926_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17569_ net758 _01857_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14323__464 clknet_1_0__leaf__08465_ VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__inv_2
XFILLER_0_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13961__246 clknet_1_1__leaf__08356_ VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__inv_2
XFILLER_0_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14033__310 clknet_1_0__leaf__08364_ VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__inv_2
X_09825_ net2151 _05402_ _05474_ VGND VGND VPWR VPWR _05484_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09756_ _05441_ _05281_ _05442_ _05275_ _05444_ VGND VGND VPWR VPWR _05445_ sky130_fd_sc_hd__o221a_1
X_12764__214 clknet_1_1__leaf__07224_ VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__inv_2
X_08707_ _04404_ _04425_ _04426_ VGND VGND VPWR VPWR _04427_ sky130_fd_sc_hd__o21a_1
X_09687_ _04916_ _05375_ _05377_ _04974_ _05378_ VGND VGND VPWR VPWR _05379_ sky130_fd_sc_hd__o221a_1
XFILLER_0_96_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_87_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14406__539 clknet_1_1__leaf__02656_ VGND VGND VPWR VPWR net571 sky130_fd_sc_hd__inv_2
X_08638_ CPU.aluIn1\[27\] _04229_ VGND VGND VPWR VPWR _04358_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_120_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08569_ CPU.aluIn1\[2\] _04288_ VGND VGND VPWR VPWR _04289_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_25_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10600_ net1414 _05968_ _05982_ _05980_ VGND VGND VPWR VPWR _02188_ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11580_ _06512_ _05911_ VGND VGND VPWR VPWR _06525_ sky130_fd_sc_hd__nor2_2
X_14298__441 clknet_1_0__leaf__08463_ VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__inv_2
XFILLER_0_18_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10531_ net1402 _05892_ _05933_ _05885_ VGND VGND VPWR VPWR _02208_ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13250_ CPU.registerFile\[19\]\[10\] _07383_ _07682_ VGND VGND VPWR VPWR _07683_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_135_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10462_ _04553_ _04555_ _04556_ VGND VGND VPWR VPWR _05875_ sky130_fd_sc_hd__and3_1
XFILLER_0_150_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12201_ net2479 _06884_ _06862_ VGND VGND VPWR VPWR _06885_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13181_ _07380_ _07611_ _07615_ _07584_ VGND VGND VPWR VPWR _07616_ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10393_ _05821_ _05822_ VGND VGND VPWR VPWR _05823_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12132_ _06838_ VGND VGND VPWR VPWR _01509_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16940_ net235 _01266_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_12063_ _05130_ net1849 _06794_ VGND VGND VPWR VPWR _06802_ sky130_fd_sc_hd__mux2_1
X_14190__369 clknet_1_0__leaf__08428_ VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__inv_2
X_14764__861 clknet_1_0__leaf__02692_ VGND VGND VPWR VPWR net893 sky130_fd_sc_hd__inv_2
X_11014_ _06209_ VGND VGND VPWR VPWR _02002_ sky130_fd_sc_hd__clkbuf_1
X_16871_ per_uart.uart0.rx_count16\[0\] _04153_ per_uart.uart0.rx_count16\[1\] VGND
+ VGND VPWR VPWR _04157_ sky130_fd_sc_hd__a21oi_1
X_16524__191 clknet_1_1__leaf__03964_ VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__inv_2
X_15822_ CPU.registerFile\[28\]\[12\] _02791_ VGND VGND VPWR VPWR _03309_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_51_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15753_ CPU.registerFile\[8\]\[10\] CPU.registerFile\[12\]\[10\] _02999_ VGND VGND
+ VPWR VPWR _03242_ sky130_fd_sc_hd__mux2_1
X_12965_ CPU.registerFile\[31\]\[2\] _07403_ _07404_ CPU.registerFile\[27\]\[2\] _07405_
+ VGND VGND VPWR VPWR _07406_ sky130_fd_sc_hd__o221a_1
X_11916_ _06724_ VGND VGND VPWR VPWR _01612_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15684_ _02797_ _03172_ _03173_ _03174_ _03054_ VGND VGND VPWR VPWR _03175_ sky130_fd_sc_hd__a221o_1
X_12896_ _07273_ _07336_ _07337_ VGND VGND VPWR VPWR _07338_ sky130_fd_sc_hd__o21a_1
XANTENNA_340 _03079_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_351 _05381_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_362 _07657_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17423_ net612 _01711_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[16\] sky130_fd_sc_hd__dfxtp_1
X_11847_ CPU.registerFile\[10\]\[20\] _05694_ _06686_ VGND VGND VPWR VPWR _06688_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_373 _07256_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_384 _05541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_395 _08014_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17354_ net543 _01642_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_11778_ _06651_ VGND VGND VPWR VPWR _01677_ sky130_fd_sc_hd__clkbuf_1
X_13517_ CPU.registerFile\[8\]\[18\] CPU.registerFile\[12\]\[18\] _07315_ VGND VGND
+ VPWR VPWR _07942_ sky130_fd_sc_hd__mux2_1
X_16305_ _03771_ _03777_ _02879_ VGND VGND VPWR VPWR _03778_ sky130_fd_sc_hd__o21a_1
X_17285_ net474 _01573_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_10729_ _06058_ VGND VGND VPWR VPWR _02136_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16236_ CPU.registerFile\[27\]\[24\] CPU.registerFile\[31\]\[24\] _08403_ VGND VGND
+ VPWR VPWR _03711_ sky130_fd_sc_hd__mux2_1
X_13448_ _07873_ _07874_ _07785_ VGND VGND VPWR VPWR _07875_ sky130_fd_sc_hd__mux2_1
Xclkload12 clknet_leaf_15_clk VGND VGND VPWR VPWR clkload12/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_151_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload23 clknet_leaf_6_clk VGND VGND VPWR VPWR clkload23/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_153_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload34 clknet_1_0__leaf__02751_ VGND VGND VPWR VPWR clkload34/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload45 clknet_1_1__leaf__02721_ VGND VGND VPWR VPWR clkload45/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload56 clknet_1_0__leaf__02699_ VGND VGND VPWR VPWR clkload56/Y sky130_fd_sc_hd__clkinvlp_4
X_16167_ _02858_ _03641_ _03643_ _02864_ VGND VGND VPWR VPWR _03644_ sky130_fd_sc_hd__a211o_1
XFILLER_0_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13379_ CPU.registerFile\[5\]\[14\] _07804_ _07807_ _07368_ VGND VGND VPWR VPWR _07808_
+ sky130_fd_sc_hd__o211a_1
Xclkload67 clknet_1_0__leaf__02682_ VGND VGND VPWR VPWR clkload67/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_50_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload78 clknet_1_0__leaf__02666_ VGND VGND VPWR VPWR clkload78/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload89 clknet_1_0__leaf__02655_ VGND VGND VPWR VPWR clkload89/Y sky130_fd_sc_hd__clkinvlp_4
X_14847__936 clknet_1_0__leaf__02700_ VGND VGND VPWR VPWR net968 sky130_fd_sc_hd__inv_2
XFILLER_0_62_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16098_ _02901_ _03575_ _03576_ _03030_ VGND VGND VPWR VPWR _03577_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_71_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_10_Left_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09610_ _05287_ _05295_ _05304_ VGND VGND VPWR VPWR _05305_ sky130_fd_sc_hd__or3_4
X_09541_ _04860_ _04886_ VGND VGND VPWR VPWR _05238_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_69_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09472_ mapped_spi_ram.rcv_data\[19\] _04688_ _04709_ mapped_spi_flash.rcv_data\[19\]
+ VGND VGND VPWR VPWR _05172_ sky130_fd_sc_hd__a22oi_4
XTAP_TAPCELL_ROW_102_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14893__978 clknet_1_1__leaf__02704_ VGND VGND VPWR VPWR net1010 sky130_fd_sc_hd__inv_2
XFILLER_0_18_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_82_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload6 clknet_leaf_27_clk VGND VGND VPWR VPWR clkload6/Y sky130_fd_sc_hd__inv_6
XFILLER_0_41_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_89_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09808_ _05475_ VGND VGND VPWR VPWR _02521_ sky130_fd_sc_hd__clkbuf_1
X_09739_ CPU.aluIn1\[0\] _04302_ VGND VGND VPWR VPWR _05428_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11701_ mapped_spi_ram.rcv_data\[10\] _06603_ _06604_ _06594_ VGND VGND VPWR VPWR
+ _01706_ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12681_ CPU.cycles\[25\] _07166_ net1428 VGND VGND VPWR VPWR _07169_ sky130_fd_sc_hd__a21oi_1
X_11632_ mapped_spi_ram.snd_bitcount\[3\] _06549_ VGND VGND VPWR VPWR _06560_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14351_ clknet_1_0__leaf__08433_ VGND VGND VPWR VPWR _08468_ sky130_fd_sc_hd__buf_1
XFILLER_0_107_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11563_ _06493_ VGND VGND VPWR VPWR _06512_ sky130_fd_sc_hd__buf_2
XFILLER_0_52_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14986__1061 clknet_1_0__leaf__02714_ VGND VGND VPWR VPWR net1093 sky130_fd_sc_hd__inv_2
X_13302_ CPU.registerFile\[9\]\[11\] _07363_ _07733_ VGND VGND VPWR VPWR _07734_ sky130_fd_sc_hd__o21a_1
X_17070_ net328 _01392_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_10514_ _05886_ _05919_ VGND VGND VPWR VPWR _05920_ sky130_fd_sc_hd__nor2_1
X_14282_ CPU.PC\[1\] _08456_ VGND VGND VPWR VPWR _08461_ sky130_fd_sc_hd__or2b_1
XFILLER_0_122_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11494_ _06464_ VGND VGND VPWR VPWR _01777_ sky130_fd_sc_hd__clkbuf_1
X_14005__286 clknet_1_1__leaf__08360_ VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_133_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16021_ CPU.registerFile\[15\]\[18\] CPU.registerFile\[11\]\[18\] _02906_ VGND VGND
+ VPWR VPWR _03502_ sky130_fd_sc_hd__mux2_1
X_13233_ CPU.registerFile\[13\]\[9\] _07629_ _07488_ CPU.registerFile\[9\]\[9\] _07489_
+ VGND VGND VPWR VPWR _07667_ sky130_fd_sc_hd__o221a_1
X_10445_ net1360 _05850_ _05851_ _05861_ VGND VGND VPWR VPWR _05862_ sky130_fd_sc_hd__a211o_1
X_13164_ _07411_ _07596_ _07599_ VGND VGND VPWR VPWR _07600_ sky130_fd_sc_hd__or3_2
XFILLER_0_20_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__02690_ _02690_ VGND VGND VPWR VPWR clknet_0__02690_ sky130_fd_sc_hd__clkbuf_16
X_10376_ _05553_ net2494 _05776_ VGND VGND VPWR VPWR _05810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12115_ _06829_ VGND VGND VPWR VPWR _01517_ sky130_fd_sc_hd__clkbuf_1
X_13095_ CPU.mem_wdata\[5\] _07229_ _07532_ _07135_ VGND VGND VPWR VPWR _01300_ sky130_fd_sc_hd__o211a_1
X_17972_ net1160 _02256_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_14352__490 clknet_1_1__leaf__08468_ VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__inv_2
X_12046_ _04958_ net2040 _06783_ VGND VGND VPWR VPWR _06793_ sky130_fd_sc_hd__mux2_1
X_16923_ CPU.mem_wdata\[7\] _04180_ _04190_ _05844_ VGND VGND VPWR VPWR _02645_ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13990__272 clknet_1_1__leaf__08359_ VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_148_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16854_ net1592 VGND VGND VPWR VPWR _02621_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_148_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15805_ CPU.registerFile\[22\]\[11\] CPU.registerFile\[23\]\[11\] _02828_ VGND VGND
+ VPWR VPWR _03293_ sky130_fd_sc_hd__mux2_1
X_16785_ _05288_ _04039_ _04975_ VGND VGND VPWR VPWR _04097_ sky130_fd_sc_hd__a21o_1
XFILLER_0_153_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_834 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15736_ CPU.registerFile\[5\]\[10\] CPU.registerFile\[4\]\[10\] _02898_ VGND VGND
+ VPWR VPWR _03225_ sky130_fd_sc_hd__mux2_1
X_12948_ CPU.registerFile\[4\]\[2\] _07388_ VGND VGND VPWR VPWR _07389_ sky130_fd_sc_hd__or2_1
X_12879_ _07316_ _07319_ _07320_ VGND VGND VPWR VPWR _07321_ sky130_fd_sc_hd__mux2_1
XANTENNA_170 _07404_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15667_ CPU.aluIn1\[7\] _03081_ _03158_ _03080_ VGND VGND VPWR VPWR _02421_ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_181 _07555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_192 _07841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_134_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17406_ net595 _01694_ VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dfxtp_2
X_14618_ clknet_1_0__leaf__02675_ VGND VGND VPWR VPWR _02678_ sky130_fd_sc_hd__buf_1
X_15598_ _03086_ _03090_ _02784_ VGND VGND VPWR VPWR _03091_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_64_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17337_ net526 _01625_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload101 clknet_1_1__leaf__08365_ VGND VGND VPWR VPWR clkload101/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_71_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17268_ net458 _01556_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[29\] sky130_fd_sc_hd__dfxtp_1
Xclkload112 clknet_1_0__leaf__03989_ VGND VGND VPWR VPWR clkload112/Y sky130_fd_sc_hd__clkinvlp_4
Xclkbuf_1_1__f__08433_ clknet_0__08433_ VGND VGND VPWR VPWR clknet_1_1__leaf__08433_
+ sky130_fd_sc_hd__clkbuf_16
X_16219_ _02856_ _03692_ _03694_ _02965_ VGND VGND VPWR VPWR _03695_ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17199_ clknet_leaf_11_clk _01487_ VGND VGND VPWR VPWR CPU.Bimm\[9\] sky130_fd_sc_hd__dfxtp_2
X_14435__565 clknet_1_0__leaf__02659_ VGND VGND VPWR VPWR net597 sky130_fd_sc_hd__inv_2
Xclkbuf_0__08464_ _08464_ VGND VGND VPWR VPWR clknet_0__08464_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__08364_ clknet_0__08364_ VGND VGND VPWR VPWR clknet_1_1__leaf__08364_
+ sky130_fd_sc_hd__clkbuf_16
X_08972_ _04690_ VGND VGND VPWR VPWR _04691_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09524_ _04317_ _04214_ _04219_ CPU.aluReg\[9\] _05221_ VGND VGND VPWR VPWR _05222_
+ sky130_fd_sc_hd__a221o_1
X_14901__985 clknet_1_0__leaf__02705_ VGND VGND VPWR VPWR net1017 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_84_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600__713 clknet_1_1__leaf__02676_ VGND VGND VPWR VPWR net745 sky130_fd_sc_hd__inv_2
X_09455_ _04955_ _05155_ _04208_ _04498_ VGND VGND VPWR VPWR _05156_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_94_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09386_ CPU.registerFile\[16\]\[16\] _05090_ _04983_ VGND VGND VPWR VPWR _05091_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_814 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14256__428 clknet_1_0__leaf__08435_ VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_115_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10230_ net1985 _05729_ _05713_ VGND VGND VPWR VPWR _05730_ sky130_fd_sc_hd__mux2_1
X_10161_ _04779_ VGND VGND VPWR VPWR _05683_ sky130_fd_sc_hd__buf_2
X_10092_ net1723 _04958_ _05633_ VGND VGND VPWR VPWR _05643_ sky130_fd_sc_hd__mux2_1
X_13920_ CPU.registerFile\[18\]\[31\] CPU.registerFile\[22\]\[31\] _07457_ VGND VGND
+ VPWR VPWR _08332_ sky130_fd_sc_hd__mux2_1
X_13851_ net1517 _08018_ _08265_ _08017_ VGND VGND VPWR VPWR _01323_ sky130_fd_sc_hd__o211a_1
X_12802_ _05337_ VGND VGND VPWR VPWR _07245_ sky130_fd_sc_hd__clkbuf_4
X_13782_ CPU.registerFile\[9\]\[26\] _07619_ _08198_ VGND VGND VPWR VPWR _08199_ sky130_fd_sc_hd__o21a_1
X_10994_ net2260 _05708_ _06190_ VGND VGND VPWR VPWR _06199_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14876__962 clknet_1_0__leaf__02703_ VGND VGND VPWR VPWR net994 sky130_fd_sc_hd__inv_2
X_15521_ CPU.registerFile\[27\]\[4\] CPU.registerFile\[31\]\[4\] _02852_ VGND VGND
+ VPWR VPWR _03016_ sky130_fd_sc_hd__mux2_1
X_12733_ _07211_ net1676 _07205_ VGND VGND VPWR VPWR _07212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15452_ _02948_ VGND VGND VPWR VPWR _02949_ sky130_fd_sc_hd__buf_4
X_18240_ net81 _02520_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_12664_ _07158_ _07159_ VGND VGND VPWR VPWR _00024_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11615_ net1387 _06494_ _06546_ _06539_ VGND VGND VPWR VPWR _01734_ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18171_ net202 _02451_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_15383_ _02772_ VGND VGND VPWR VPWR _02881_ sky130_fd_sc_hd__buf_4
XFILLER_0_143_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12595_ CPU.mem_wbusy _06865_ _07120_ VGND VGND VPWR VPWR _07121_ sky130_fd_sc_hd__or3b_1
XFILLER_0_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17122_ clknet_leaf_17_clk _00024_ VGND VGND VPWR VPWR CPU.cycles\[18\] sky130_fd_sc_hd__dfxtp_1
X_11546_ net1409 _06499_ _06489_ VGND VGND VPWR VPWR _06500_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17053_ net311 _01375_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_14265_ _04802_ _04947_ _04962_ _08443_ VGND VGND VPWR VPWR _08444_ sky130_fd_sc_hd__or4_1
Xclkbuf_1_1__f__02711_ clknet_0__02711_ VGND VGND VPWR VPWR clknet_1_1__leaf__02711_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11477_ _05532_ CPU.registerFile\[25\]\[11\] _06455_ VGND VGND VPWR VPWR _06456_
+ sky130_fd_sc_hd__mux2_1
X_16004_ _02924_ _03483_ _03484_ _03485_ _02782_ VGND VGND VPWR VPWR _03486_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13216_ _07417_ VGND VGND VPWR VPWR _07650_ sky130_fd_sc_hd__buf_4
XFILLER_0_111_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10428_ _05848_ VGND VGND VPWR VPWR _02226_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13147_ _07369_ _07580_ _07582_ _07392_ VGND VGND VPWR VPWR _07583_ sky130_fd_sc_hd__a211o_1
Xclkbuf_0__02673_ _02673_ VGND VGND VPWR VPWR clknet_0__02673_ sky130_fd_sc_hd__clkbuf_16
X_10359_ _05801_ VGND VGND VPWR VPWR _02249_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13078_ CPU.registerFile\[14\]\[5\] CPU.registerFile\[10\]\[5\] _07274_ VGND VGND
+ VPWR VPWR _07516_ sky130_fd_sc_hd__mux2_1
X_17955_ net1143 _02239_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_12029_ _06784_ VGND VGND VPWR VPWR _01558_ sky130_fd_sc_hd__clkbuf_1
X_16906_ _04616_ _04615_ _04612_ _04640_ VGND VGND VPWR VPWR _04181_ sky130_fd_sc_hd__and4_1
X_17886_ net1075 _02170_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[4\] sky130_fd_sc_hd__dfxtp_1
X_16837_ per_uart.uart0.txd_reg\[7\] per_uart.d_in_uart\[7\] _07178_ VGND VGND VPWR
+ VPWR _04135_ sky130_fd_sc_hd__mux2_1
X_16768_ _04052_ _05043_ _08453_ VGND VGND VPWR VPWR _04083_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_66_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15719_ CPU.registerFile\[30\]\[9\] CPU.registerFile\[26\]\[9\] _02881_ VGND VGND
+ VPWR VPWR _03209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16699_ _08457_ _04022_ _04023_ _04024_ VGND VGND VPWR VPWR _04025_ sky130_fd_sc_hd__a31o_1
X_16587__59 clknet_1_0__leaf__03969_ VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__inv_2
X_09240_ CPU.PC\[22\] _04821_ VGND VGND VPWR VPWR _04951_ sky130_fd_sc_hd__xor2_1
XFILLER_0_7_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09171_ _04864_ _04882_ _04862_ VGND VGND VPWR VPWR _04883_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_32_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18369_ net37 _02647_ VGND VGND VPWR VPWR mapped_spi_ram.div_counter\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_32_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_778 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__03989_ _03989_ VGND VGND VPWR VPWR clknet_0__03989_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_98_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_131_Right_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08955_ _04478_ _04673_ VGND VGND VPWR VPWR _04674_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_102_Left_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08886_ _04566_ _04605_ _04565_ VGND VGND VPWR VPWR _04606_ sky130_fd_sc_hd__a21oi_1
X_14985__1060 clknet_1_0__leaf__02714_ VGND VGND VPWR VPWR net1092 sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__02662_ clknet_0__02662_ VGND VGND VPWR VPWR clknet_1_0__leaf__02662_
+ sky130_fd_sc_hd__clkbuf_16
X_09507_ _05199_ _05205_ _04492_ VGND VGND VPWR VPWR _05206_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_67_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09438_ _04504_ _04812_ _04503_ CPU.cycles\[13\] _05139_ VGND VGND VPWR VPWR _05140_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_111_Left_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09369_ CPU.aluIn1\[16\] _04254_ _04699_ VGND VGND VPWR VPWR _05074_ sky130_fd_sc_hd__o21a_1
XFILLER_0_136_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11400_ _05524_ net2190 _06408_ VGND VGND VPWR VPWR _06415_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12380_ _07007_ VGND VGND VPWR VPWR _01396_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_70 _05108_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_81 _05208_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11331_ _05524_ net2138 _06371_ VGND VGND VPWR VPWR _06378_ sky130_fd_sc_hd__mux2_1
XANTENNA_92 _05306_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11262_ _06341_ VGND VGND VPWR VPWR _01886_ sky130_fd_sc_hd__clkbuf_1
X_13001_ _07232_ _07433_ _07440_ VGND VGND VPWR VPWR _07441_ sky130_fd_sc_hd__a21o_1
X_10213_ _05718_ VGND VGND VPWR VPWR _02327_ sky130_fd_sc_hd__clkbuf_1
X_11193_ _05522_ net1778 _06299_ VGND VGND VPWR VPWR _06305_ sky130_fd_sc_hd__mux2_1
X_10144_ net2011 _05668_ _05671_ VGND VGND VPWR VPWR _05672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17740_ net929 _02024_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_128_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10075_ _05634_ VGND VGND VPWR VPWR _02381_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_128_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13903_ CPU.registerFile\[30\]\[30\] CPU.registerFile\[26\]\[30\] _07297_ VGND VGND
+ VPWR VPWR _08316_ sky130_fd_sc_hd__mux2_1
X_17671_ net860 _01959_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_16622_ _03986_ VGND VGND VPWR VPWR _02548_ sky130_fd_sc_hd__clkbuf_1
X_13834_ _08241_ _08248_ _07411_ VGND VGND VPWR VPWR _08249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14464__591 clknet_1_0__leaf__02662_ VGND VGND VPWR VPWR net623 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_141_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13765_ CPU.registerFile\[18\]\[26\] CPU.registerFile\[22\]\[26\] _07315_ VGND VGND
+ VPWR VPWR _08182_ sky130_fd_sc_hd__mux2_1
X_10977_ _06178_ VGND VGND VPWR VPWR _06190_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_0__f__08367_ clknet_0__08367_ VGND VGND VPWR VPWR clknet_1_0__leaf__08367_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_84_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15504_ _02851_ VGND VGND VPWR VPWR _02999_ sky130_fd_sc_hd__clkbuf_8
X_12716_ _07195_ _07196_ _07197_ VGND VGND VPWR VPWR _07198_ sky130_fd_sc_hd__or3_1
XFILLER_0_84_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13696_ _07801_ _08112_ _08113_ _08114_ _07555_ VGND VGND VPWR VPWR _08115_ sky130_fd_sc_hd__a221o_1
X_16484_ CPU.registerFile\[25\]\[31\] CPU.registerFile\[29\]\[31\] _03254_ VGND VGND
+ VPWR VPWR _03952_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18223_ net64 _02503_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12647_ _07148_ _07149_ VGND VGND VPWR VPWR _00017_ sky130_fd_sc_hd__nor2_1
X_15435_ _02922_ _02931_ _02879_ VGND VGND VPWR VPWR _02932_ sky130_fd_sc_hd__a21o_1
XFILLER_0_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15366_ _08396_ VGND VGND VPWR VPWR _02864_ sky130_fd_sc_hd__buf_4
X_18154_ clknet_leaf_26_clk _02434_ VGND VGND VPWR VPWR CPU.aluIn1\[20\] sky130_fd_sc_hd__dfxtp_4
X_12578_ _07112_ VGND VGND VPWR VPWR _01270_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14239__412 clknet_1_1__leaf__08434_ VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__inv_2
XFILLER_0_81_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17105_ clknet_leaf_23_clk _00026_ VGND VGND VPWR VPWR CPU.cycles\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11529_ _06490_ VGND VGND VPWR VPWR _06491_ sky130_fd_sc_hd__inv_2
X_18085_ net148 _02365_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_15297_ _02769_ VGND VGND VPWR VPWR _02796_ sky130_fd_sc_hd__buf_4
XFILLER_0_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold307 CPU.rs2\[14\] VGND VGND VPWR VPWR net1548 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold318 CPU.registerFile\[16\]\[19\] VGND VGND VPWR VPWR net1559 sky130_fd_sc_hd__dlygate4sd3_1
Xhold329 CPU.registerFile\[5\]\[28\] VGND VGND VPWR VPWR net1570 sky130_fd_sc_hd__dlygate4sd3_1
X_17036_ net294 _01358_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14179_ _08427_ VGND VGND VPWR VPWR _01489_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14950__1029 clknet_1_0__leaf__02710_ VGND VGND VPWR VPWR net1061 sky130_fd_sc_hd__inv_2
Xclkbuf_0__02656_ _02656_ VGND VGND VPWR VPWR clknet_0__02656_ sky130_fd_sc_hd__clkbuf_16
X_08740_ CPU.aluIn1\[23\] _04237_ VGND VGND VPWR VPWR _04460_ sky130_fd_sc_hd__nand2_1
Xhold1007 CPU.registerFile\[30\]\[19\] VGND VGND VPWR VPWR net2248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1018 CPU.registerFile\[7\]\[16\] VGND VGND VPWR VPWR net2259 sky130_fd_sc_hd__dlygate4sd3_1
X_17938_ net1127 _02222_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[18\] sky130_fd_sc_hd__dfxtp_1
Xhold1029 CPU.aluReg\[0\] VGND VGND VPWR VPWR net2270 sky130_fd_sc_hd__dlygate4sd3_1
X_14547__666 clknet_1_1__leaf__02670_ VGND VGND VPWR VPWR net698 sky130_fd_sc_hd__inv_2
X_08671_ CPU.aluIn1\[15\] VGND VGND VPWR VPWR _04391_ sky130_fd_sc_hd__inv_2
X_17869_ net1058 _02153_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[27\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_37_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09223_ _04934_ VGND VGND VPWR VPWR _02573_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_840 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_756 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09154_ _04499_ CPU.Iimm\[4\] _04665_ _04830_ VGND VGND VPWR VPWR _04866_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14712__814 clknet_1_0__leaf__02687_ VGND VGND VPWR VPWR net846 sky130_fd_sc_hd__inv_2
XFILLER_0_71_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09085_ _04797_ VGND VGND VPWR VPWR _04798_ sky130_fd_sc_hd__clkbuf_4
X_14292__436 clknet_1_0__leaf__08462_ VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__inv_2
XFILLER_0_130_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold830 CPU.registerFile\[26\]\[5\] VGND VGND VPWR VPWR net2071 sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 CPU.registerFile\[19\]\[3\] VGND VGND VPWR VPWR net2082 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold852 CPU.registerFile\[1\]\[30\] VGND VGND VPWR VPWR net2093 sky130_fd_sc_hd__dlygate4sd3_1
Xhold863 CPU.registerFile\[2\]\[22\] VGND VGND VPWR VPWR net2104 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold874 CPU.PC\[2\] VGND VGND VPWR VPWR net2115 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold885 CPU.registerFile\[22\]\[1\] VGND VGND VPWR VPWR net2126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 CPU.registerFile\[13\]\[1\] VGND VGND VPWR VPWR net2137 sky130_fd_sc_hd__dlygate4sd3_1
X_09987_ _05586_ VGND VGND VPWR VPWR _02453_ sky130_fd_sc_hd__clkbuf_1
X_08938_ _04493_ _04657_ VGND VGND VPWR VPWR _04658_ sky130_fd_sc_hd__or2_2
X_08869_ _04505_ VGND VGND VPWR VPWR _04589_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_98_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10900_ _06149_ VGND VGND VPWR VPWR _02056_ sky130_fd_sc_hd__clkbuf_1
X_11880_ net2521 _05727_ _06697_ VGND VGND VPWR VPWR _06705_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__02714_ clknet_0__02714_ VGND VGND VPWR VPWR clknet_1_0__leaf__02714_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_123_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10831_ _06112_ VGND VGND VPWR VPWR _02088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_123_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13550_ CPU.registerFile\[15\]\[19\] _07482_ _07973_ _07621_ _07483_ VGND VGND VPWR
+ VPWR _07974_ sky130_fd_sc_hd__o221a_1
XFILLER_0_67_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10762_ _05501_ net1693 _06070_ VGND VGND VPWR VPWR _06076_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12501_ net1913 _05712_ _07071_ VGND VGND VPWR VPWR _07072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13481_ _07584_ _07896_ _07899_ _07906_ VGND VGND VPWR VPWR _07907_ sky130_fd_sc_hd__o31a_1
XFILLER_0_82_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10693_ _06039_ VGND VGND VPWR VPWR _02153_ sky130_fd_sc_hd__clkbuf_1
X_12432_ _07012_ VGND VGND VPWR VPWR _07035_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_152_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12363_ _06998_ VGND VGND VPWR VPWR _01404_ sky130_fd_sc_hd__clkbuf_1
X_14102_ _04499_ VGND VGND VPWR VPWR _08379_ sky130_fd_sc_hd__clkbuf_2
X_11314_ _05507_ net2159 _06360_ VGND VGND VPWR VPWR _06369_ sky130_fd_sc_hd__mux2_1
X_15082_ _07180_ _02725_ _02727_ VGND VGND VPWR VPWR _02271_ sky130_fd_sc_hd__a21oi_1
X_12294_ CPU.aluIn1\[6\] _06955_ _06927_ VGND VGND VPWR VPWR _06956_ sky130_fd_sc_hd__mux2_1
X_11245_ _06332_ VGND VGND VPWR VPWR _01894_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11176_ _05505_ net1767 _06288_ VGND VGND VPWR VPWR _06296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10127_ _05661_ VGND VGND VPWR VPWR _02356_ sky130_fd_sc_hd__clkbuf_1
X_15984_ CPU.registerFile\[6\]\[17\] _02819_ VGND VGND VPWR VPWR _03466_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_143_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17723_ net912 _02007_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_10058_ _05624_ VGND VGND VPWR VPWR _02388_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17654_ net843 _01942_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_16605_ per_uart.uart0.rx_bitcount\[3\] per_uart.uart0.rx_bitcount\[2\] per_uart.uart0.rx_bitcount\[1\]
+ per_uart.uart0.rx_bitcount\[0\] VGND VGND VPWR VPWR _03976_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_34_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13817_ _07334_ _08222_ _08225_ _08232_ _07766_ VGND VGND VPWR VPWR _08233_ sky130_fd_sc_hd__o311a_1
X_17585_ net774 _01873_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13748_ CPU.registerFile\[2\]\[25\] CPU.registerFile\[10\]\[25\] _07304_ VGND VGND
+ VPWR VPWR _08166_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_158_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_158_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16467_ CPU.registerFile\[22\]\[31\] _08399_ VGND VGND VPWR VPWR _03935_ sky130_fd_sc_hd__and2_1
X_13679_ _07639_ _08096_ _08097_ _08098_ _07570_ VGND VGND VPWR VPWR _08099_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18206_ net47 _02486_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15418_ CPU.registerFile\[9\]\[2\] CPU.registerFile\[13\]\[2\] _02887_ VGND VGND
+ VPWR VPWR _02915_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16398_ _03864_ _03867_ _02858_ VGND VGND VPWR VPWR _03868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18137_ clknet_leaf_27_clk _02417_ VGND VGND VPWR VPWR CPU.aluIn1\[3\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_143_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15349_ CPU.aluIn1\[0\] _08018_ _02847_ _08017_ VGND VGND VPWR VPWR _02414_ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold104 mapped_spi_ram.cmd_addr\[23\] VGND VGND VPWR VPWR net1345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 _07141_ VGND VGND VPWR VPWR net1356 sky130_fd_sc_hd__dlygate4sd3_1
X_18068_ net1241 _02348_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[30\] sky130_fd_sc_hd__dfxtp_1
Xhold126 mapped_spi_flash.cmd_addr\[3\] VGND VGND VPWR VPWR net1367 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold137 mapped_spi_ram.cmd_addr\[13\] VGND VGND VPWR VPWR net1378 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold148 mapped_spi_ram.cmd_addr\[20\] VGND VGND VPWR VPWR net1389 sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ _05541_ net2293 _05533_ VGND VGND VPWR VPWR _05542_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17019_ net277 _01341_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[13\] sky130_fd_sc_hd__dfxtp_1
Xhold159 mapped_spi_flash.cmd_addr\[11\] VGND VGND VPWR VPWR net1400 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09841_ _04713_ VGND VGND VPWR VPWR _05495_ sky130_fd_sc_hd__buf_6
Xclkbuf_0__02708_ _02708_ VGND VGND VPWR VPWR clknet_0__02708_ sky130_fd_sc_hd__clkbuf_16
X_09772_ _05456_ VGND VGND VPWR VPWR _02538_ sky130_fd_sc_hd__clkbuf_1
X_08723_ _04390_ _04441_ _04442_ VGND VGND VPWR VPWR _04443_ sky130_fd_sc_hd__o21a_1
X_14480__606 clknet_1_0__leaf__02663_ VGND VGND VPWR VPWR net638 sky130_fd_sc_hd__inv_2
XFILLER_0_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08654_ _04373_ VGND VGND VPWR VPWR _04374_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_68_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08585_ CPU.aluIn1\[3\] _04286_ VGND VGND VPWR VPWR _04305_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_105_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09206_ CPU.PC\[5\] _04917_ VGND VGND VPWR VPWR _04918_ sky130_fd_sc_hd__and2_1
XFILLER_0_147_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14300__443 clknet_1_0__leaf__08463_ VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__inv_2
XFILLER_0_51_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09137_ CPU.PC\[13\] _04847_ VGND VGND VPWR VPWR _04849_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_20_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09068_ _04781_ VGND VGND VPWR VPWR _02575_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold660 CPU.registerFile\[29\]\[8\] VGND VGND VPWR VPWR net1901 sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 CPU.registerFile\[7\]\[9\] VGND VGND VPWR VPWR net1912 sky130_fd_sc_hd__dlygate4sd3_1
X_11030_ _06218_ VGND VGND VPWR VPWR _01995_ sky130_fd_sc_hd__clkbuf_1
Xhold682 CPU.registerFile\[19\]\[19\] VGND VGND VPWR VPWR net1923 sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 per_uart.d_in_uart\[5\] VGND VGND VPWR VPWR net1934 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_125_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12981_ _07418_ _07419_ _07421_ VGND VGND VPWR VPWR _07422_ sky130_fd_sc_hd__o21a_1
X_11932_ _06732_ VGND VGND VPWR VPWR _01604_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11863_ net2418 _05710_ _06686_ VGND VGND VPWR VPWR _06696_ sky130_fd_sc_hd__mux2_1
X_14651_ clknet_1_0__leaf__02675_ VGND VGND VPWR VPWR _02681_ sky130_fd_sc_hd__buf_1
XFILLER_0_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13602_ CPU.registerFile\[15\]\[21\] _07772_ _07773_ CPU.registerFile\[11\]\[21\]
+ _08023_ VGND VGND VPWR VPWR _08024_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_28_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10814_ _05553_ net1781 _06069_ VGND VGND VPWR VPWR _06103_ sky130_fd_sc_hd__mux2_1
X_17370_ net559 _01658_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11794_ _06659_ VGND VGND VPWR VPWR _01669_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16321_ _05384_ _03790_ _03793_ VGND VGND VPWR VPWR _03794_ sky130_fd_sc_hd__or3_1
XFILLER_0_27_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10745_ _06066_ VGND VGND VPWR VPWR _02128_ sky130_fd_sc_hd__clkbuf_1
X_13533_ CPU.registerFile\[16\]\[19\] CPU.registerFile\[20\]\[19\] _07233_ VGND VGND
+ VPWR VPWR _07957_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13464_ _07475_ _07889_ _07890_ VGND VGND VPWR VPWR _07891_ sky130_fd_sc_hd__o21a_1
X_16252_ _02926_ _03725_ _03726_ VGND VGND VPWR VPWR _03727_ sky130_fd_sc_hd__o21a_1
X_10676_ _06022_ _06018_ mapped_spi_flash.rcv_bitcount\[0\] VGND VGND VPWR VPWR _06029_
+ sky130_fd_sc_hd__mux2_1
X_14576__692 clknet_1_0__leaf__02673_ VGND VGND VPWR VPWR net724 sky130_fd_sc_hd__inv_2
X_12415_ _07026_ VGND VGND VPWR VPWR _01380_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13395_ CPU.registerFile\[13\]\[14\] _07361_ _07521_ CPU.registerFile\[9\]\[14\]
+ _07285_ VGND VGND VPWR VPWR _07824_ sky130_fd_sc_hd__o221a_1
X_16183_ CPU.registerFile\[2\]\[22\] _03143_ _02822_ CPU.registerFile\[3\]\[22\] _03144_
+ VGND VGND VPWR VPWR _03660_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_136_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_153_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12346_ _05008_ net2086 _06988_ VGND VGND VPWR VPWR _06990_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12277_ CPU.aluReg\[11\] CPU.aluReg\[9\] _06939_ VGND VGND VPWR VPWR _06943_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11228_ _05594_ _06250_ VGND VGND VPWR VPWR _06323_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_56_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11159_ _06286_ VGND VGND VPWR VPWR _01934_ sky130_fd_sc_hd__clkbuf_1
X_15967_ CPU.registerFile\[6\]\[16\] _03057_ _03140_ _03449_ VGND VGND VPWR VPWR _03450_
+ sky130_fd_sc_hd__o211a_1
X_14741__840 clknet_1_0__leaf__02690_ VGND VGND VPWR VPWR net872 sky130_fd_sc_hd__inv_2
X_17706_ net895 _01994_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_15898_ _03378_ _03382_ _03138_ VGND VGND VPWR VPWR _03383_ sky130_fd_sc_hd__a21o_1
X_16501__170 clknet_1_1__leaf__03962_ VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__inv_2
X_17637_ net826 _01925_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17568_ net757 _01856_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14659__767 clknet_1_1__leaf__02681_ VGND VGND VPWR VPWR net799 sky130_fd_sc_hd__inv_2
XFILLER_0_147_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17499_ net688 _01787_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14824__915 clknet_1_1__leaf__02698_ VGND VGND VPWR VPWR net947 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_6_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09824_ _05483_ VGND VGND VPWR VPWR _02513_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_107_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09755_ mapped_spi_ram.rcv_data\[24\] _04783_ _05277_ _05443_ VGND VGND VPWR VPWR
+ _05444_ sky130_fd_sc_hd__a211o_1
X_08706_ _04315_ _04271_ VGND VGND VPWR VPWR _04426_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09686_ CPU.cycles\[3\] _04502_ VGND VGND VPWR VPWR _05378_ sky130_fd_sc_hd__nand2_1
X_08637_ _04354_ _04234_ _04356_ VGND VGND VPWR VPWR _04357_ sky130_fd_sc_hd__a21oi_2
XTAP_TAPCELL_ROW_87_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08568_ CPU.mem_wdata\[2\] CPU.Iimm\[2\] _04202_ VGND VGND VPWR VPWR _04288_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_25_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08499_ _04218_ VGND VGND VPWR VPWR _04219_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14870__957 clknet_1_1__leaf__02702_ VGND VGND VPWR VPWR net989 sky130_fd_sc_hd__inv_2
X_10530_ net1367 _05887_ _05856_ _05932_ VGND VGND VPWR VPWR _05933_ sky130_fd_sc_hd__a211o_1
XFILLER_0_146_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10461_ net1399 _05849_ _05874_ _05855_ VGND VGND VPWR VPWR _02219_ sky130_fd_sc_hd__o211a_1
X_12200_ CPU.aluIn1\[28\] _06883_ _06865_ VGND VGND VPWR VPWR _06884_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_118_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13180_ _07369_ _07612_ _07614_ _07392_ VGND VGND VPWR VPWR _07615_ sky130_fd_sc_hd__a211o_1
X_10392_ CPU.mem_rstrb _04784_ _05812_ VGND VGND VPWR VPWR _05822_ sky130_fd_sc_hd__a21oi_1
X_12131_ _05130_ net1751 _06830_ VGND VGND VPWR VPWR _06838_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12062_ _06801_ VGND VGND VPWR VPWR _01542_ sky130_fd_sc_hd__clkbuf_1
Xhold490 CPU.registerFile\[22\]\[31\] VGND VGND VPWR VPWR net1731 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11013_ net1563 _05727_ _06201_ VGND VGND VPWR VPWR _06209_ sky130_fd_sc_hd__mux2_1
X_16870_ per_uart.uart0.rx_count16\[1\] per_uart.uart0.rx_count16\[0\] _04153_ VGND
+ VGND VPWR VPWR _04156_ sky130_fd_sc_hd__and3_1
X_15821_ CPU.registerFile\[30\]\[12\] CPU.registerFile\[26\]\[12\] _02787_ VGND VGND
+ VPWR VPWR _03308_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_51_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15752_ _08411_ _03232_ _03240_ _02935_ VGND VGND VPWR VPWR _03241_ sky130_fd_sc_hd__o211a_1
X_12964_ _07252_ VGND VGND VPWR VPWR _07405_ sky130_fd_sc_hd__clkbuf_8
Xhold1190 CPU.registerFile\[8\]\[8\] VGND VGND VPWR VPWR net2431 sky130_fd_sc_hd__dlygate4sd3_1
X_11915_ CPU.registerFile\[11\]\[20\] _05694_ _06722_ VGND VGND VPWR VPWR _06724_
+ sky130_fd_sc_hd__mux2_1
X_15683_ CPU.registerFile\[25\]\[8\] _02802_ _02803_ VGND VGND VPWR VPWR _03174_ sky130_fd_sc_hd__o21a_1
X_12895_ CPU.registerFile\[15\]\[1\] _07276_ _07277_ CPU.registerFile\[11\]\[1\] _07278_
+ VGND VGND VPWR VPWR _07337_ sky130_fd_sc_hd__o221a_1
XFILLER_0_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_330 CPU.mem_wdata\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_341 _05050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_352 _05511_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17422_ net611 _01710_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[15\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_363 _02806_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11846_ _06687_ VGND VGND VPWR VPWR _01645_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_374 _07277_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_385 _05541_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_396 _02786_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17353_ net542 _01641_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[17\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_138_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ _04982_ net1928 _06650_ VGND VGND VPWR VPWR _06651_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16304_ _08401_ _03773_ _03776_ _02844_ VGND VGND VPWR VPWR _03777_ sky130_fd_sc_hd__o211a_1
X_13516_ _07412_ _07939_ _07940_ VGND VGND VPWR VPWR _07941_ sky130_fd_sc_hd__o21a_1
X_10728_ _05535_ CPU.registerFile\[28\]\[10\] _06056_ VGND VGND VPWR VPWR _06058_
+ sky130_fd_sc_hd__mux2_1
X_17284_ net473 _01572_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14496_ clknet_1_1__leaf__02664_ VGND VGND VPWR VPWR _02666_ sky130_fd_sc_hd__buf_1
XFILLER_0_83_798 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_153_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16235_ _02911_ _03707_ _03709_ _03245_ VGND VGND VPWR VPWR _03710_ sky130_fd_sc_hd__a211o_1
XFILLER_0_152_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13447_ CPU.registerFile\[6\]\[16\] CPU.registerFile\[7\]\[16\] _07311_ VGND VGND
+ VPWR VPWR _07874_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_889 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10659_ _05820_ _06015_ _06016_ VGND VGND VPWR VPWR _06017_ sky130_fd_sc_hd__a21oi_1
Xclkload13 clknet_leaf_16_clk VGND VGND VPWR VPWR clkload13/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload24 clknet_leaf_8_clk VGND VGND VPWR VPWR clkload24/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_58_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload35 clknet_1_1__leaf__02750_ VGND VGND VPWR VPWR clkload35/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload46 clknet_1_0__leaf__02708_ VGND VGND VPWR VPWR clkload46/X sky130_fd_sc_hd__clkbuf_8
X_13378_ CPU.registerFile\[4\]\[14\] _07374_ VGND VGND VPWR VPWR _07807_ sky130_fd_sc_hd__or2_1
X_16166_ CPU.registerFile\[24\]\[22\] _02816_ _05071_ _03642_ VGND VGND VPWR VPWR
+ _03643_ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload57 clknet_1_1__leaf__02698_ VGND VGND VPWR VPWR clkload57/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload68 clknet_1_0__leaf__02681_ VGND VGND VPWR VPWR clkload68/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload79 clknet_1_0__leaf__02665_ VGND VGND VPWR VPWR clkload79/Y sky130_fd_sc_hd__clkinvlp_4
X_12329_ _04731_ net1788 _06977_ VGND VGND VPWR VPWR _06981_ sky130_fd_sc_hd__mux2_1
X_16097_ CPU.registerFile\[19\]\[20\] CPU.registerFile\[17\]\[20\] _03025_ VGND VGND
+ VPWR VPWR _03576_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16999_ clknet_leaf_21_clk _01325_ VGND VGND VPWR VPWR CPU.rs2\[30\] sky130_fd_sc_hd__dfxtp_1
X_09540_ _04716_ _05236_ _04717_ VGND VGND VPWR VPWR _05237_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09471_ _05171_ VGND VGND VPWR VPWR _02562_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_69_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14592__707 clknet_1_1__leaf__02674_ VGND VGND VPWR VPWR net739 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_82_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload7 clknet_leaf_28_clk VGND VGND VPWR VPWR clkload7/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_132_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16657__2 clknet_1_0__leaf__07220_ VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__inv_2
XFILLER_0_15_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14412__544 clknet_1_1__leaf__02657_ VGND VGND VPWR VPWR net576 sky130_fd_sc_hd__inv_2
XFILLER_0_100_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09807_ net1990 _05188_ _05474_ VGND VGND VPWR VPWR _05475_ sky130_fd_sc_hd__mux2_1
X_09738_ _05427_ VGND VGND VPWR VPWR _02551_ sky130_fd_sc_hd__clkbuf_1
X_09669_ mapped_spi_ram.rcv_data\[11\] _04783_ _04784_ mapped_spi_flash.rcv_data\[11\]
+ VGND VGND VPWR VPWR _05361_ sky130_fd_sc_hd__a22o_4
X_11700_ mapped_spi_ram.rcv_data\[11\] _06601_ VGND VGND VPWR VPWR _06604_ sky130_fd_sc_hd__or2_1
X_12680_ CPU.cycles\[25\] CPU.cycles\[26\] _07166_ VGND VGND VPWR VPWR _07168_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11631_ net1474 _06555_ _06559_ _06474_ VGND VGND VPWR VPWR _01731_ sky130_fd_sc_hd__o22a_1
XFILLER_0_126_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11562_ net1390 _06495_ _06511_ _06006_ VGND VGND VPWR VPWR _01752_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_145_Right_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13301_ CPU.registerFile\[13\]\[11\] _07402_ _07732_ _07621_ _07249_ VGND VGND VPWR
+ VPWR _07733_ sky130_fd_sc_hd__o221a_1
XFILLER_0_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10513_ CPU.PC\[7\] _05867_ _05917_ _05918_ VGND VGND VPWR VPWR _05919_ sky130_fd_sc_hd__o2bb2a_1
X_14281_ _08436_ _08459_ _05412_ VGND VGND VPWR VPWR _08460_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11493_ _05549_ net2371 _06455_ VGND VGND VPWR VPWR _06464_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13232_ CPU.registerFile\[8\]\[9\] CPU.registerFile\[12\]\[9\] _07265_ VGND VGND
+ VPWR VPWR _07666_ sky130_fd_sc_hd__mux2_1
X_16020_ _02786_ _03498_ _03500_ _03019_ VGND VGND VPWR VPWR _03501_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_133_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10444_ _05852_ _04611_ VGND VGND VPWR VPWR _05861_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13163_ _07475_ _07597_ _07598_ VGND VGND VPWR VPWR _07599_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10375_ _05809_ VGND VGND VPWR VPWR _02241_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12114_ _04958_ net1997 _06819_ VGND VGND VPWR VPWR _06829_ sky130_fd_sc_hd__mux2_1
X_13094_ _07230_ _07515_ _07531_ _07309_ VGND VGND VPWR VPWR _07532_ sky130_fd_sc_hd__a211o_1
X_17971_ net1159 _02255_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_14688__793 clknet_1_0__leaf__02684_ VGND VGND VPWR VPWR net825 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_53_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12045_ _06792_ VGND VGND VPWR VPWR _01550_ sky130_fd_sc_hd__clkbuf_1
X_16922_ net1747 _04182_ VGND VGND VPWR VPWR _04190_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14387__521 clknet_1_1__leaf__02655_ VGND VGND VPWR VPWR net553 sky130_fd_sc_hd__inv_2
XFILLER_0_137_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16853_ net1591 per_uart.rx_data\[5\] _04139_ VGND VGND VPWR VPWR _04145_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_148_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15804_ _03065_ _03290_ _03291_ VGND VGND VPWR VPWR _03292_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16784_ _04032_ net2481 VGND VGND VPWR VPWR _04096_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_148_Left_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15735_ CPU.aluIn1\[9\] _02958_ _03207_ _03224_ _02995_ VGND VGND VPWR VPWR _02423_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_88_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12947_ _05337_ VGND VGND VPWR VPWR _07388_ sky130_fd_sc_hd__buf_4
XFILLER_0_87_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14086__359 clknet_1_1__leaf__08368_ VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__inv_2
XFILLER_0_158_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15666_ _02757_ _03128_ _03139_ _03157_ _02846_ VGND VGND VPWR VPWR _03158_ sky130_fd_sc_hd__a311o_2
X_12878_ _04971_ VGND VGND VPWR VPWR _07320_ sky130_fd_sc_hd__buf_8
XANTENNA_160 _07320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_171 _07412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_182 _07555_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17405_ net594 _01693_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_bitcount\[5\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_193 _07841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11829_ _06678_ VGND VGND VPWR VPWR _01653_ sky130_fd_sc_hd__clkbuf_1
X_15597_ _02771_ _03087_ _03088_ _03089_ _02782_ VGND VGND VPWR VPWR _03090_ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14853__941 clknet_1_0__leaf__02701_ VGND VGND VPWR VPWR net973 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_16_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17336_ net525 _01624_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_112_Right_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17267_ net457 _01555_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[28\] sky130_fd_sc_hd__dfxtp_1
Xclkload102 clknet_1_1__leaf__08364_ VGND VGND VPWR VPWR clkload102/Y sky130_fd_sc_hd__clkinvlp_4
XPHY_EDGE_ROW_157_Left_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload113 clknet_1_0__leaf__03970_ VGND VGND VPWR VPWR clkload113/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_71_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16218_ _02796_ _03693_ VGND VGND VPWR VPWR _03694_ sky130_fd_sc_hd__or2_1
Xclkbuf_1_1__f__08432_ clknet_0__08432_ VGND VGND VPWR VPWR clknet_1_1__leaf__08432_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17198_ clknet_leaf_11_clk _01486_ VGND VGND VPWR VPWR CPU.Bimm\[8\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_11_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_470 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__08463_ _08463_ VGND VGND VPWR VPWR clknet_0__08463_ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f__08363_ clknet_0__08363_ VGND VGND VPWR VPWR clknet_1_1__leaf__08363_
+ sky130_fd_sc_hd__clkbuf_16
X_16149_ CPU.registerFile\[18\]\[21\] _03068_ _03069_ CPU.registerFile\[19\]\[21\]
+ _03074_ VGND VGND VPWR VPWR _03627_ sky130_fd_sc_hd__o221a_1
XFILLER_0_141_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08971_ _04618_ VGND VGND VPWR VPWR _04690_ sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09523_ _04428_ _04701_ _04210_ _04269_ VGND VGND VPWR VPWR _05221_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_149_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09454_ CPU.PC\[12\] _04922_ VGND VGND VPWR VPWR _05155_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09385_ _05089_ VGND VGND VPWR VPWR _05090_ sky130_fd_sc_hd__buf_6
XFILLER_0_143_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10160_ _05682_ VGND VGND VPWR VPWR _02344_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10091_ _05642_ VGND VGND VPWR VPWR _02373_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13850_ _07397_ _08249_ _08264_ _08015_ VGND VGND VPWR VPWR _08265_ sky130_fd_sc_hd__a211o_1
XFILLER_0_16_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15237__146 clknet_1_0__leaf__02754_ VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__inv_2
X_12801_ _07235_ VGND VGND VPWR VPWR _07244_ sky130_fd_sc_hd__buf_4
X_13781_ CPU.registerFile\[13\]\[26\] _07629_ _08197_ _07371_ _04971_ VGND VGND VPWR
+ VPWR _08198_ sky130_fd_sc_hd__o221a_1
X_10993_ _06198_ VGND VGND VPWR VPWR _02012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15520_ _02764_ VGND VGND VPWR VPWR _03015_ sky130_fd_sc_hd__buf_4
X_14011__291 clknet_1_1__leaf__08361_ VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__inv_2
X_12732_ per_uart.d_in_uart\[3\] _07178_ _07203_ per_uart.uart0.txd_reg\[4\] VGND
+ VGND VPWR VPWR _07211_ sky130_fd_sc_hd__a22o_1
X_15451_ _05010_ VGND VGND VPWR VPWR _02948_ sky130_fd_sc_hd__buf_4
XFILLER_0_155_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12663_ net1411 _07156_ VGND VGND VPWR VPWR _07159_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18170_ net201 _02450_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_11614_ net1930 _06501_ _06496_ CPU.mem_wdata\[1\] _06508_ VGND VGND VPWR VPWR _06546_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15382_ _02866_ _02878_ _02879_ VGND VGND VPWR VPWR _02880_ sky130_fd_sc_hd__o21a_1
XFILLER_0_154_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12594_ mapped_spi_flash.rbusy mapped_spi_ram.rbusy VGND VGND VPWR VPWR _07120_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17121_ clknet_leaf_17_clk _00023_ VGND VGND VPWR VPWR CPU.cycles\[17\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11545_ _06493_ VGND VGND VPWR VPWR _06499_ sky130_fd_sc_hd__buf_2
XFILLER_0_135_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17052_ net310 _01374_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[14\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__02710_ clknet_0__02710_ VGND VGND VPWR VPWR clknet_1_1__leaf__02710_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_40_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14264_ _04997_ _05014_ _05037_ _08442_ VGND VGND VPWR VPWR _08443_ sky130_fd_sc_hd__or4_1
X_11476_ _06432_ VGND VGND VPWR VPWR _06455_ sky130_fd_sc_hd__clkbuf_4
X_16003_ CPU.registerFile\[13\]\[17\] _02775_ VGND VGND VPWR VPWR _03485_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10427_ _05830_ _05847_ VGND VGND VPWR VPWR _05848_ sky130_fd_sc_hd__and2_1
X_13215_ CPU.registerFile\[18\]\[9\] CPU.registerFile\[22\]\[9\] _07648_ VGND VGND
+ VPWR VPWR _07649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13146_ CPU.registerFile\[3\]\[7\] _04987_ _07581_ _04939_ VGND VGND VPWR VPWR _07582_
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_0__02672_ _02672_ VGND VGND VPWR VPWR clknet_0__02672_ sky130_fd_sc_hd__clkbuf_16
X_10358_ _05535_ net2462 _05799_ VGND VGND VPWR VPWR _05801_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13077_ _07507_ _07513_ _07514_ VGND VGND VPWR VPWR _07515_ sky130_fd_sc_hd__mux2_1
X_17954_ net1142 _02238_ VGND VGND VPWR VPWR mapped_spi_flash.rbusy sky130_fd_sc_hd__dfxtp_1
X_10289_ _05535_ CPU.registerFile\[20\]\[10\] _05762_ VGND VGND VPWR VPWR _05764_
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12028_ _04659_ net1642 _06783_ VGND VGND VPWR VPWR _06784_ sky130_fd_sc_hd__mux2_1
X_16905_ net1290 _06468_ VGND VGND VPWR VPWR _04180_ sky130_fd_sc_hd__nand2_2
X_17885_ net1074 _02169_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[3\] sky130_fd_sc_hd__dfxtp_1
X_16836_ net2296 _04126_ _04134_ _04115_ VGND VGND VPWR VPWR _02614_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16767_ _04027_ _04039_ _05042_ VGND VGND VPWR VPWR _04082_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_66_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15718_ CPU.registerFile\[28\]\[9\] CPU.registerFile\[24\]\[9\] _02881_ VGND VGND
+ VPWR VPWR _03208_ sky130_fd_sc_hd__mux2_1
X_16698_ _04001_ _05263_ _03990_ VGND VGND VPWR VPWR _04024_ sky130_fd_sc_hd__a21o_1
XFILLER_0_158_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15649_ CPU.registerFile\[7\]\[7\] _05092_ VGND VGND VPWR VPWR _03141_ sky130_fd_sc_hd__or2_1
X_14441__570 clknet_1_1__leaf__02660_ VGND VGND VPWR VPWR net602 sky130_fd_sc_hd__inv_2
XFILLER_0_118_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09170_ _04865_ _04880_ _04881_ VGND VGND VPWR VPWR _04882_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18368_ net36 _02646_ VGND VGND VPWR VPWR mapped_spi_ram.div_counter\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_32_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17319_ net508 _01607_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18299_ net33 _02579_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14359__497 clknet_1_0__leaf__08468_ VGND VGND VPWR VPWR net529 sky130_fd_sc_hd__inv_2
XFILLER_0_114_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__03988_ _03988_ VGND VGND VPWR VPWR clknet_0__03988_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_52_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13997__279 clknet_1_0__leaf__08359_ VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__inv_2
XFILLER_0_11_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08954_ _04378_ _04477_ _04367_ VGND VGND VPWR VPWR _04673_ sky130_fd_sc_hd__or3b_1
X_08885_ _04564_ _04569_ _04568_ VGND VGND VPWR VPWR _04605_ sky130_fd_sc_hd__a21o_1
X_14069__343 clknet_1_1__leaf__08367_ VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__inv_2
X_14524__645 clknet_1_0__leaf__02668_ VGND VGND VPWR VPWR net677 sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__02661_ clknet_0__02661_ VGND VGND VPWR VPWR clknet_1_0__leaf__02661_
+ sky130_fd_sc_hd__clkbuf_16
X_09506_ _04267_ _04489_ _05204_ _04679_ VGND VGND VPWR VPWR _05205_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09437_ _04817_ _05136_ _05138_ _04915_ VGND VGND VPWR VPWR _05139_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_137_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15027__1099 clknet_1_1__leaf__02717_ VGND VGND VPWR VPWR net1131 sky130_fd_sc_hd__inv_2
XFILLER_0_19_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09368_ CPU.Jimm\[16\] _04812_ _04989_ CPU.cycles\[16\] VGND VGND VPWR VPWR _05073_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09299_ _05007_ VGND VGND VPWR VPWR _05008_ sky130_fd_sc_hd__buf_6
XFILLER_0_151_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_60 _05046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_71 _05108_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_82 _05229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11330_ _06377_ VGND VGND VPWR VPWR _01854_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_97_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_93 _05306_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11261_ CPU.registerFile\[9\]\[16\] _05702_ _06335_ VGND VGND VPWR VPWR _06341_ sky130_fd_sc_hd__mux2_1
X_14570__687 clknet_1_0__leaf__02672_ VGND VGND VPWR VPWR net719 sky130_fd_sc_hd__inv_2
XFILLER_0_30_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13000_ _07254_ _07435_ _07439_ _07268_ VGND VGND VPWR VPWR _07440_ sky130_fd_sc_hd__o211a_1
X_10212_ net1909 _05717_ _05713_ VGND VGND VPWR VPWR _05718_ sky130_fd_sc_hd__mux2_1
X_11192_ _06304_ VGND VGND VPWR VPWR _01919_ sky130_fd_sc_hd__clkbuf_1
X_10143_ _05670_ VGND VGND VPWR VPWR _05671_ sky130_fd_sc_hd__buf_4
X_10074_ net2007 _04659_ _05633_ VGND VGND VPWR VPWR _05634_ sky130_fd_sc_hd__mux2_1
X_14951_ clknet_1_0__leaf__02708_ VGND VGND VPWR VPWR _02711_ sky130_fd_sc_hd__buf_1
XFILLER_0_27_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13902_ _07519_ _08313_ _08314_ VGND VGND VPWR VPWR _08315_ sky130_fd_sc_hd__o21a_1
X_17670_ net859 _01958_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_16621_ net1825 net1797 _03979_ VGND VGND VPWR VPWR _03986_ sky130_fd_sc_hd__mux2_1
X_13833_ _08244_ _08247_ _07253_ VGND VGND VPWR VPWR _08248_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__08435_ clknet_0__08435_ VGND VGND VPWR VPWR clknet_1_0__leaf__08435_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_18_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13764_ _07254_ _08176_ _08180_ _07646_ VGND VGND VPWR VPWR _08181_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_48_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14499__622 clknet_1_0__leaf__02666_ VGND VGND VPWR VPWR net654 sky130_fd_sc_hd__inv_2
X_10976_ _06189_ VGND VGND VPWR VPWR _02020_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__08366_ clknet_0__08366_ VGND VGND VPWR VPWR clknet_1_0__leaf__08366_
+ sky130_fd_sc_hd__clkbuf_16
X_15503_ _02996_ _02997_ _02856_ VGND VGND VPWR VPWR _02998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12715_ per_uart.uart0.tx_count16\[3\] per_uart.uart0.tx_count16\[2\] per_uart.tx_busy
+ VGND VGND VPWR VPWR _07197_ sky130_fd_sc_hd__or3b_1
X_16483_ _03946_ _03950_ _02784_ VGND VGND VPWR VPWR _03951_ sky130_fd_sc_hd__a21o_1
X_13695_ CPU.registerFile\[3\]\[24\] _07804_ _07987_ VGND VGND VPWR VPWR _08114_ sky130_fd_sc_hd__o21a_1
X_18222_ net63 _02502_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15434_ _02924_ _02925_ _02927_ _02929_ _02930_ VGND VGND VPWR VPWR _02931_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_61_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12646_ CPU.cycles\[10\] _07146_ net1403 VGND VGND VPWR VPWR _07149_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18153_ clknet_leaf_28_clk _02433_ VGND VGND VPWR VPWR CPU.aluIn1\[19\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_143_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15365_ CPU.registerFile\[12\]\[1\] _02826_ _02860_ _02862_ VGND VGND VPWR VPWR _02863_
+ sky130_fd_sc_hd__o211a_1
X_12577_ net1636 _05272_ _07107_ VGND VGND VPWR VPWR _07112_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16592__63 clknet_1_1__leaf__03970_ VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__inv_2
X_17104_ clknet_leaf_24_clk _00015_ VGND VGND VPWR VPWR CPU.cycles\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18084_ net147 _02364_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_11528_ mapped_spi_ram.state\[1\] _06487_ VGND VGND VPWR VPWR _06490_ sky130_fd_sc_hd__and2_1
XFILLER_0_151_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15296_ _02786_ _02788_ _02793_ _02794_ VGND VGND VPWR VPWR _02795_ sky130_fd_sc_hd__a211o_1
XFILLER_0_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold308 CPU.PC\[5\] VGND VGND VPWR VPWR net1549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold319 CPU.registerFile\[14\]\[1\] VGND VGND VPWR VPWR net1560 sky130_fd_sc_hd__dlygate4sd3_1
X_17035_ net293 _01357_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_14247_ clknet_1_1__leaf__08433_ VGND VGND VPWR VPWR _08435_ sky130_fd_sc_hd__buf_1
X_11459_ _06446_ VGND VGND VPWR VPWR _01794_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__02724_ _02724_ VGND VGND VPWR VPWR clknet_0__02724_ sky130_fd_sc_hd__clkbuf_16
X_14178_ _04496_ _08426_ _07127_ VGND VGND VPWR VPWR _08427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0__02655_ _02655_ VGND VGND VPWR VPWR clknet_0__02655_ sky130_fd_sc_hd__clkbuf_16
X_13129_ _07230_ _07547_ _07565_ _07309_ VGND VGND VPWR VPWR _07566_ sky130_fd_sc_hd__a211o_1
Xhold1008 CPU.registerFile\[10\]\[31\] VGND VGND VPWR VPWR net2249 sky130_fd_sc_hd__dlygate4sd3_1
X_15059__1125 clknet_1_0__leaf__02722_ VGND VGND VPWR VPWR net1157 sky130_fd_sc_hd__inv_2
X_17937_ net1126 _02221_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[17\] sky130_fd_sc_hd__dfxtp_1
Xhold1019 CPU.registerFile\[6\]\[13\] VGND VGND VPWR VPWR net2260 sky130_fd_sc_hd__dlygate4sd3_1
X_08670_ _04389_ _04254_ VGND VGND VPWR VPWR _04390_ sky130_fd_sc_hd__nor2_1
X_17868_ net1057 _02152_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_16819_ net1546 _04121_ _04122_ _03632_ VGND VGND VPWR VPWR _02609_ sky130_fd_sc_hd__o211a_1
X_17799_ net988 _02083_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[21\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_37_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09222_ net1687 _04933_ _04668_ VGND VGND VPWR VPWR _04934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09153_ CPU.Bimm\[5\] _04819_ CPU.PC\[5\] VGND VGND VPWR VPWR _04865_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09084_ CPU.cycles\[24\] _04687_ _04786_ _04796_ VGND VGND VPWR VPWR _04797_ sky130_fd_sc_hd__a211o_2
XTAP_TAPCELL_ROW_79_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold820 CPU.registerFile\[3\]\[5\] VGND VGND VPWR VPWR net2061 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold831 CPU.registerFile\[21\]\[27\] VGND VGND VPWR VPWR net2072 sky130_fd_sc_hd__dlygate4sd3_1
Xhold842 CPU.registerFile\[26\]\[23\] VGND VGND VPWR VPWR net2083 sky130_fd_sc_hd__dlygate4sd3_1
X_15151__1179 clknet_1_0__leaf__02745_ VGND VGND VPWR VPWR net1211 sky130_fd_sc_hd__inv_2
Xhold853 CPU.registerFile\[7\]\[13\] VGND VGND VPWR VPWR net2094 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_782 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold864 CPU.registerFile\[19\]\[12\] VGND VGND VPWR VPWR net2105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 CPU.registerFile\[7\]\[14\] VGND VGND VPWR VPWR net2116 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_92_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold886 CPU.registerFile\[26\]\[28\] VGND VGND VPWR VPWR net2127 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__08429_ _08429_ VGND VGND VPWR VPWR clknet_0__08429_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold897 CPU.registerFile\[23\]\[15\] VGND VGND VPWR VPWR net2138 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09986_ _05541_ net2088 _05581_ VGND VGND VPWR VPWR _05586_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08937_ _04496_ _04498_ _04503_ CPU.cycles\[31\] _04656_ VGND VGND VPWR VPWR _04657_
+ sky130_fd_sc_hd__a221o_1
X_08868_ _04506_ _04584_ _04585_ _04587_ VGND VGND VPWR VPWR _04588_ sky130_fd_sc_hd__o31a_2
Xclkbuf_1_0__f__02713_ clknet_0__02713_ VGND VGND VPWR VPWR clknet_1_0__leaf__02713_
+ sky130_fd_sc_hd__clkbuf_16
X_08799_ CPU.aluIn1\[4\] _04517_ VGND VGND VPWR VPWR _04519_ sky130_fd_sc_hd__or2_1
X_10830_ net1663 _05681_ _06106_ VGND VGND VPWR VPWR _06112_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_123_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10761_ _06075_ VGND VGND VPWR VPWR _02121_ sky130_fd_sc_hd__clkbuf_1
X_12500_ _07048_ VGND VGND VPWR VPWR _07071_ sky130_fd_sc_hd__clkbuf_4
X_13480_ _07271_ _07902_ _07905_ _07306_ VGND VGND VPWR VPWR _07906_ sky130_fd_sc_hd__o31a_1
X_10692_ _05499_ net1721 _06034_ VGND VGND VPWR VPWR _06039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12431_ _07034_ VGND VGND VPWR VPWR _01372_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12362_ _05170_ net1734 _06988_ VGND VGND VPWR VPWR _06998_ sky130_fd_sc_hd__mux2_1
X_14101_ _08378_ VGND VGND VPWR VPWR _01460_ sky130_fd_sc_hd__clkbuf_1
X_11313_ _06368_ VGND VGND VPWR VPWR _01862_ sky130_fd_sc_hd__clkbuf_1
X_15081_ _02726_ VGND VGND VPWR VPWR _02727_ sky130_fd_sc_hd__buf_2
X_12293_ CPU.aluReg\[7\] CPU.aluReg\[5\] _06939_ VGND VGND VPWR VPWR _06955_ sky130_fd_sc_hd__mux2_1
X_11244_ net1897 _05685_ _06324_ VGND VGND VPWR VPWR _06332_ sky130_fd_sc_hd__mux2_1
X_14032_ clknet_1_0__leaf__08363_ VGND VGND VPWR VPWR _08364_ sky130_fd_sc_hd__buf_1
XFILLER_0_31_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11175_ _06295_ VGND VGND VPWR VPWR _01927_ sky130_fd_sc_hd__clkbuf_1
X_10126_ net1910 _05306_ _05655_ VGND VGND VPWR VPWR _05661_ sky130_fd_sc_hd__mux2_1
X_15983_ CPU.registerFile\[1\]\[17\] _03030_ _03464_ _03028_ VGND VGND VPWR VPWR _03465_
+ sky130_fd_sc_hd__a22o_1
X_16629__75 clknet_1_0__leaf__03971_ VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__inv_2
X_17722_ net911 _02006_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_10057_ net1921 _05306_ _05618_ VGND VGND VPWR VPWR _05624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17653_ net842 _01941_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_16644__89 clknet_1_0__leaf__03988_ VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__inv_2
X_16604_ per_uart.uart0.rx_bitcount\[2\] per_uart.uart0.rx_bitcount\[1\] per_uart.uart0.rx_bitcount\[0\]
+ per_uart.uart0.rx_bitcount\[3\] VGND VGND VPWR VPWR _03975_ sky130_fd_sc_hd__and4bb_1
X_13816_ _07405_ _08228_ _08229_ _08231_ _07359_ VGND VGND VPWR VPWR _08232_ sky130_fd_sc_hd__a221o_1
X_17584_ net773 _01872_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13747_ _07474_ _08161_ _08164_ VGND VGND VPWR VPWR _08165_ sky130_fd_sc_hd__or3_1
X_10959_ net1611 _05673_ _06179_ VGND VGND VPWR VPWR _06181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_668 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_158_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_158_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16466_ CPU.registerFile\[21\]\[31\] CPU.registerFile\[23\]\[31\] _02769_ VGND VGND
+ VPWR VPWR _03934_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_158_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13678_ CPU.registerFile\[2\]\[23\] _07417_ _07376_ VGND VGND VPWR VPWR _08098_ sky130_fd_sc_hd__o21a_1
XFILLER_0_6_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18205_ net46 _02485_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_15417_ _05071_ VGND VGND VPWR VPWR _02914_ sky130_fd_sc_hd__buf_4
X_12629_ _07138_ _07139_ VGND VGND VPWR VPWR _00040_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16397_ CPU.registerFile\[2\]\[29\] _03227_ _03228_ CPU.registerFile\[3\]\[29\] _03866_
+ VGND VGND VPWR VPWR _03867_ sky130_fd_sc_hd__a221o_1
X_18136_ clknet_leaf_27_clk _02416_ VGND VGND VPWR VPWR CPU.aluIn1\[2\] sky130_fd_sc_hd__dfxtp_4
X_15348_ _02757_ _02785_ _02811_ _02845_ _02846_ VGND VGND VPWR VPWR _02847_ sky130_fd_sc_hd__a311o_2
XPHY_EDGE_ROW_130_Left_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18067_ net1240 _02347_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_14553__671 clknet_1_1__leaf__02671_ VGND VGND VPWR VPWR net703 sky130_fd_sc_hd__inv_2
Xhold105 mapped_spi_flash.rcv_bitcount\[3\] VGND VGND VPWR VPWR net1346 sky130_fd_sc_hd__dlygate4sd3_1
X_15279_ _02777_ VGND VGND VPWR VPWR _02778_ sky130_fd_sc_hd__clkbuf_4
Xhold116 mapped_spi_flash.rcv_bitcount\[2\] VGND VGND VPWR VPWR net1357 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 mapped_spi_flash.cmd_addr\[14\] VGND VGND VPWR VPWR net1368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 CPU.cycles\[20\] VGND VGND VPWR VPWR net1379 sky130_fd_sc_hd__dlygate4sd3_1
X_17018_ net276 _01340_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[12\] sky130_fd_sc_hd__dfxtp_1
Xhold149 mapped_spi_ram.cmd_addr\[19\] VGND VGND VPWR VPWR net1390 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__02707_ _02707_ VGND VGND VPWR VPWR clknet_0__02707_ sky130_fd_sc_hd__clkbuf_16
X_09840_ _05494_ VGND VGND VPWR VPWR _02508_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15026__1098 clknet_1_1__leaf__02717_ VGND VGND VPWR VPWR net1130 sky130_fd_sc_hd__inv_2
X_09771_ net1803 _04731_ _05452_ VGND VGND VPWR VPWR _05456_ sky130_fd_sc_hd__mux2_1
X_08722_ _04253_ _04252_ VGND VGND VPWR VPWR _04442_ sky130_fd_sc_hd__nand2_2
X_08653_ CPU.Bimm\[10\] _04372_ VGND VGND VPWR VPWR _04373_ sky130_fd_sc_hd__and2_2
XFILLER_0_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_922 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08584_ _04300_ _04302_ CPU.aluIn1\[0\] _04303_ VGND VGND VPWR VPWR _04304_ sky130_fd_sc_hd__a31oi_4
XTAP_TAPCELL_ROW_105_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16556__30 clknet_1_0__leaf__03967_ VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__inv_2
XFILLER_0_45_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09205_ CPU.PC\[4\] CPU.PC\[3\] CPU.PC\[2\] VGND VGND VPWR VPWR _04917_ sky130_fd_sc_hd__and3_1
X_14636__746 clknet_1_0__leaf__02679_ VGND VGND VPWR VPWR net778 sky130_fd_sc_hd__inv_2
XFILLER_0_91_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09136_ CPU.PC\[13\] _04847_ VGND VGND VPWR VPWR _04848_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_20_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16571__44 clknet_1_0__leaf__03968_ VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__inv_2
XFILLER_0_114_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09067_ net1752 _04780_ _04668_ VGND VGND VPWR VPWR _04781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_924 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold650 CPU.registerFile\[20\]\[0\] VGND VGND VPWR VPWR net1891 sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 CPU.registerFile\[29\]\[26\] VGND VGND VPWR VPWR net1902 sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 CPU.registerFile\[3\]\[11\] VGND VGND VPWR VPWR net1913 sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 CPU.registerFile\[26\]\[26\] VGND VGND VPWR VPWR net1924 sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 CPU.registerFile\[29\]\[6\] VGND VGND VPWR VPWR net1935 sky130_fd_sc_hd__dlygate4sd3_1
X_09969_ _05524_ net1840 _05570_ VGND VGND VPWR VPWR _05577_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_125_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12980_ CPU.registerFile\[13\]\[2\] _07402_ _07420_ CPU.registerFile\[9\]\[2\] _07249_
+ VGND VGND VPWR VPWR _07421_ sky130_fd_sc_hd__o221a_1
X_14682__788 clknet_1_0__leaf__02683_ VGND VGND VPWR VPWR net820 sky130_fd_sc_hd__inv_2
X_11931_ CPU.registerFile\[11\]\[12\] _05710_ _06722_ VGND VGND VPWR VPWR _06732_
+ sky130_fd_sc_hd__mux2_1
X_14381__516 clknet_1_1__leaf__02654_ VGND VGND VPWR VPWR net548 sky130_fd_sc_hd__inv_2
XFILLER_0_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11862_ _06695_ VGND VGND VPWR VPWR _01637_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13601_ _07370_ _08022_ VGND VGND VPWR VPWR _08023_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10813_ _06102_ VGND VGND VPWR VPWR _02096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11793_ _05150_ net1837 _06650_ VGND VGND VPWR VPWR _06659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_832 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16320_ _03030_ _03791_ _03792_ _02901_ VGND VGND VPWR VPWR _03793_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13532_ CPU.registerFile\[23\]\[19\] _07362_ _07619_ CPU.registerFile\[19\]\[19\]
+ _07955_ VGND VGND VPWR VPWR _07956_ sky130_fd_sc_hd__o221a_1
XFILLER_0_39_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10744_ _05551_ CPU.registerFile\[28\]\[2\] _06056_ VGND VGND VPWR VPWR _06066_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16251_ CPU.registerFile\[18\]\[24\] _03068_ _03069_ CPU.registerFile\[19\]\[24\]
+ _03074_ VGND VGND VPWR VPWR _03726_ sky130_fd_sc_hd__o221a_1
X_13463_ CPU.registerFile\[15\]\[16\] _07402_ _07500_ CPU.registerFile\[11\]\[16\]
+ _07327_ VGND VGND VPWR VPWR _07890_ sky130_fd_sc_hd__o221a_1
XFILLER_0_125_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10675_ net1527 _06018_ _06022_ _06028_ VGND VGND VPWR VPWR _02160_ sky130_fd_sc_hd__a22o_1
X_15058__1124 clknet_1_0__leaf__02722_ VGND VGND VPWR VPWR net1156 sky130_fd_sc_hd__inv_2
XFILLER_0_152_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12414_ _05008_ net1977 _07024_ VGND VGND VPWR VPWR _07026_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16182_ CPU.registerFile\[6\]\[22\] _03026_ _03140_ _03658_ VGND VGND VPWR VPWR _03659_
+ sky130_fd_sc_hd__o211a_1
X_13394_ CPU.registerFile\[8\]\[14\] CPU.registerFile\[12\]\[14\] _07318_ VGND VGND
+ VPWR VPWR _07823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_153_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_153_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12345_ _06989_ VGND VGND VPWR VPWR _01413_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15064_ clknet_1_1__leaf__02720_ VGND VGND VPWR VPWR _02723_ sky130_fd_sc_hd__buf_1
X_12276_ _06942_ VGND VGND VPWR VPWR _01435_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11227_ _06322_ VGND VGND VPWR VPWR _01902_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_56_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11158_ CPU.registerFile\[8\]\[0\] _05735_ _06251_ VGND VGND VPWR VPWR _06286_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10109_ net2414 _05130_ _05644_ VGND VGND VPWR VPWR _05652_ sky130_fd_sc_hd__mux2_1
X_11089_ net2114 _05735_ _06214_ VGND VGND VPWR VPWR _06249_ sky130_fd_sc_hd__mux2_1
X_15966_ CPU.registerFile\[7\]\[16\] _03317_ VGND VGND VPWR VPWR _03449_ sky130_fd_sc_hd__or2_1
X_17705_ net894 _01993_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_14917_ clknet_1_1__leaf__02697_ VGND VGND VPWR VPWR _02707_ sky130_fd_sc_hd__buf_1
X_15897_ _02885_ _03379_ _03380_ _03381_ _03054_ VGND VGND VPWR VPWR _03382_ sky130_fd_sc_hd__a221o_1
XFILLER_0_157_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17636_ net825 _01924_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15150__1178 clknet_1_1__leaf__02745_ VGND VGND VPWR VPWR net1210 sky130_fd_sc_hd__inv_2
X_17567_ net756 _01855_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_17498_ net687 _01786_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16449_ _08400_ _03915_ _03916_ _03917_ _08396_ VGND VGND VPWR VPWR _03918_ sky130_fd_sc_hd__o221a_1
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18119_ net182 _02399_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14217__393 clknet_1_1__leaf__08431_ VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__inv_2
X_09823_ net2082 _05381_ _05474_ VGND VGND VPWR VPWR _05483_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09754_ mapped_spi_flash.rcv_data\[24\] _04691_ net1290 per_uart.rx_data\[0\] VGND
+ VGND VPWR VPWR _05443_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_107_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08705_ _04405_ _04423_ _04424_ VGND VGND VPWR VPWR _04425_ sky130_fd_sc_hd__o21a_1
X_09685_ _04878_ _05376_ VGND VGND VPWR VPWR _05377_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_126_Right_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08636_ _04232_ _04355_ VGND VGND VPWR VPWR _04356_ sky130_fd_sc_hd__nand2b_2
XTAP_TAPCELL_ROW_87_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08567_ CPU.aluIn1\[3\] _04286_ VGND VGND VPWR VPWR _04287_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_25_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08498_ _04217_ VGND VGND VPWR VPWR _04218_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10460_ net1368 _05850_ _05851_ _05873_ VGND VGND VPWR VPWR _05874_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_118_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09119_ _04495_ _04830_ VGND VGND VPWR VPWR _04831_ sky130_fd_sc_hd__and2_2
XFILLER_0_122_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10391_ mapped_spi_flash.clk_div _05819_ _05820_ VGND VGND VPWR VPWR _05821_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_150_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12130_ _06837_ VGND VGND VPWR VPWR _01510_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12061_ _05109_ net1826 _06794_ VGND VGND VPWR VPWR _06801_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold480 CPU.registerFile\[28\]\[27\] VGND VGND VPWR VPWR net1721 sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 CPU.registerFile\[18\]\[0\] VGND VGND VPWR VPWR net1732 sky130_fd_sc_hd__dlygate4sd3_1
X_11012_ _06208_ VGND VGND VPWR VPWR _02003_ sky130_fd_sc_hd__clkbuf_1
X_15820_ _03302_ _03306_ _02784_ VGND VGND VPWR VPWR _03307_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_51_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15751_ _02949_ _03236_ _03239_ VGND VGND VPWR VPWR _03240_ sky130_fd_sc_hd__or3_4
X_12963_ _07238_ VGND VGND VPWR VPWR _07404_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_99_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1180 CPU.registerFile\[23\]\[4\] VGND VGND VPWR VPWR net2421 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1191 CPU.registerFile\[25\]\[29\] VGND VGND VPWR VPWR net2432 sky130_fd_sc_hd__dlygate4sd3_1
X_11914_ _06723_ VGND VGND VPWR VPWR _01613_ sky130_fd_sc_hd__clkbuf_1
X_15682_ CPU.registerFile\[29\]\[8\] _02800_ VGND VGND VPWR VPWR _03173_ sky130_fd_sc_hd__or2_1
X_12894_ CPU.registerFile\[14\]\[1\] CPU.registerFile\[10\]\[1\] _07274_ VGND VGND
+ VPWR VPWR _07336_ sky130_fd_sc_hd__mux2_1
XANTENNA_320 _07914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_331 CPU.mem_wdata\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_342 _05071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17421_ net610 _01709_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[14\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_353 _05543_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11845_ net2251 _05691_ _06686_ VGND VGND VPWR VPWR _06687_ sky130_fd_sc_hd__mux2_1
XANTENNA_364 _02889_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_375 _07285_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_142_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_386 _07233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17352_ net541 _01640_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[16\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_397 _03019_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11776_ _06638_ VGND VGND VPWR VPWR _06650_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_155_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16303_ _08405_ _03774_ _03775_ VGND VGND VPWR VPWR _03776_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13515_ CPU.registerFile\[15\]\[18\] _07414_ _07326_ CPU.registerFile\[11\]\[18\]
+ _07252_ VGND VGND VPWR VPWR _07940_ sky130_fd_sc_hd__o221a_1
X_14619__730 clknet_1_0__leaf__02678_ VGND VGND VPWR VPWR net762 sky130_fd_sc_hd__inv_2
X_17283_ net472 _01571_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_10727_ _06057_ VGND VGND VPWR VPWR _02137_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15025__1097 clknet_1_1__leaf__02717_ VGND VGND VPWR VPWR net1129 sky130_fd_sc_hd__inv_2
XFILLER_0_70_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16535__11 clknet_1_1__leaf__03965_ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__inv_2
X_16234_ CPU.registerFile\[24\]\[24\] _03130_ _02780_ _03708_ VGND VGND VPWR VPWR
+ _03709_ sky130_fd_sc_hd__o211a_1
X_13446_ CPU.registerFile\[2\]\[16\] CPU.registerFile\[3\]\[16\] _07311_ VGND VGND
+ VPWR VPWR _07873_ sky130_fd_sc_hd__mux2_1
X_10658_ mapped_spi_flash.clk_div mapped_spi_flash.state\[3\] VGND VGND VPWR VPWR
+ _06016_ sky130_fd_sc_hd__and2b_1
Xclkload14 clknet_leaf_17_clk VGND VGND VPWR VPWR clkload14/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_152_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload25 clknet_leaf_9_clk VGND VGND VPWR VPWR clkload25/Y sky130_fd_sc_hd__bufinv_16
Xclkload36 clknet_1_0__leaf__07222_ VGND VGND VPWR VPWR clkload36/X sky130_fd_sc_hd__clkbuf_8
X_16165_ CPU.registerFile\[28\]\[22\] _05049_ VGND VGND VPWR VPWR _03642_ sky130_fd_sc_hd__or2_1
X_13377_ _07801_ _07802_ _07803_ _07805_ _07555_ VGND VGND VPWR VPWR _07806_ sky130_fd_sc_hd__a221o_1
XFILLER_0_106_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload47 clknet_1_0__leaf__02718_ VGND VGND VPWR VPWR clkload47/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload58 clknet_1_1__leaf__02686_ VGND VGND VPWR VPWR clkload58/X sky130_fd_sc_hd__clkbuf_8
X_10589_ mapped_spi_flash.rcv_data\[26\] _05970_ VGND VGND VPWR VPWR _05976_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload69 clknet_1_0__leaf__02678_ VGND VGND VPWR VPWR clkload69/Y sky130_fd_sc_hd__clkinvlp_4
X_16550__25 clknet_1_0__leaf__03966_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__inv_2
X_12328_ _06980_ VGND VGND VPWR VPWR _01421_ sky130_fd_sc_hd__clkbuf_1
X_16096_ CPU.registerFile\[16\]\[20\] CPU.registerFile\[18\]\[20\] _03032_ VGND VGND
+ VPWR VPWR _03575_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12259_ _06929_ VGND VGND VPWR VPWR _01439_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_71_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14665__772 clknet_1_0__leaf__02682_ VGND VGND VPWR VPWR net804 sky130_fd_sc_hd__inv_2
X_16998_ clknet_leaf_21_clk _01324_ VGND VGND VPWR VPWR CPU.rs2\[29\] sky130_fd_sc_hd__dfxtp_1
X_15949_ CPU.registerFile\[12\]\[16\] _03118_ VGND VGND VPWR VPWR _03432_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09470_ net2469 _05170_ _04983_ VGND VGND VPWR VPWR _05171_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17619_ net808 _01907_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14063__338 clknet_1_1__leaf__08366_ VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_22_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload8 clknet_leaf_29_clk VGND VGND VPWR VPWR clkload8/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_128_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14830__920 clknet_1_0__leaf__02699_ VGND VGND VPWR VPWR net952 sky130_fd_sc_hd__inv_2
XFILLER_0_15_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14748__847 clknet_1_1__leaf__02690_ VGND VGND VPWR VPWR net879 sky130_fd_sc_hd__inv_2
XFILLER_0_2_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16508__177 clknet_1_0__leaf__03962_ VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_89_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09806_ _05451_ VGND VGND VPWR VPWR _05474_ sky130_fd_sc_hd__buf_4
XFILLER_0_157_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15057__1123 clknet_1_1__leaf__02722_ VGND VGND VPWR VPWR net1155 sky130_fd_sc_hd__inv_2
X_09737_ net1600 _05426_ _04667_ VGND VGND VPWR VPWR _05427_ sky130_fd_sc_hd__mux2_1
X_09668_ _05360_ VGND VGND VPWR VPWR _02554_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08619_ _04336_ _04252_ _04250_ _04338_ VGND VGND VPWR VPWR _04339_ sky130_fd_sc_hd__a31o_4
X_09599_ _04818_ _05293_ VGND VGND VPWR VPWR _05294_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11630_ _06555_ _06558_ VGND VGND VPWR VPWR _06559_ sky130_fd_sc_hd__nand2_1
X_14794__889 clknet_1_1__leaf__02694_ VGND VGND VPWR VPWR net921 sky130_fd_sc_hd__inv_2
XFILLER_0_108_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14493__617 clknet_1_1__leaf__02665_ VGND VGND VPWR VPWR net649 sky130_fd_sc_hd__inv_2
X_11561_ net1370 _06499_ _06509_ _06510_ VGND VGND VPWR VPWR _06511_ sky130_fd_sc_hd__a211o_1
XFILLER_0_108_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13300_ CPU.registerFile\[8\]\[11\] CPU.registerFile\[12\]\[11\] _05283_ VGND VGND
+ VPWR VPWR _07732_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10512_ _04516_ _05914_ _05916_ _04629_ VGND VGND VPWR VPWR _05918_ sky130_fd_sc_hd__a31o_1
X_14280_ _08453_ VGND VGND VPWR VPWR _08459_ sky130_fd_sc_hd__buf_2
X_11492_ _06463_ VGND VGND VPWR VPWR _01778_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13231_ _07474_ _07661_ _07664_ VGND VGND VPWR VPWR _07665_ sky130_fd_sc_hd__or3_1
X_10443_ net1343 _05849_ _05860_ _05855_ VGND VGND VPWR VPWR _02223_ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13162_ CPU.registerFile\[15\]\[7\] _07402_ _07500_ CPU.registerFile\[11\]\[7\] _07483_
+ VGND VGND VPWR VPWR _07598_ sky130_fd_sc_hd__o221a_1
XFILLER_0_60_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10374_ _05551_ net1916 _05799_ VGND VGND VPWR VPWR _05809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12113_ _06828_ VGND VGND VPWR VPWR _01518_ sky130_fd_sc_hd__clkbuf_1
X_14233__408 clknet_1_1__leaf__08432_ VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__inv_2
XFILLER_0_131_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13093_ _07271_ _07518_ _07523_ _07530_ _07306_ VGND VGND VPWR VPWR _07531_ sky130_fd_sc_hd__o311a_1
X_17970_ net1158 _02254_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_53_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14807__900 clknet_1_1__leaf__02696_ VGND VGND VPWR VPWR net932 sky130_fd_sc_hd__inv_2
X_12044_ _04933_ net2083 _06783_ VGND VGND VPWR VPWR _06792_ sky130_fd_sc_hd__mux2_1
X_16921_ CPU.mem_wdata\[6\] _04180_ _04189_ _04176_ VGND VGND VPWR VPWR _02644_ sky130_fd_sc_hd__o211a_1
X_16852_ net1566 VGND VGND VPWR VPWR _02620_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_148_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747__200 clknet_1_0__leaf__07221_ VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__inv_2
X_15803_ CPU.registerFile\[16\]\[11\] _03068_ _03069_ CPU.registerFile\[17\]\[11\]
+ _02779_ VGND VGND VPWR VPWR _03291_ sky130_fd_sc_hd__o221a_1
X_16783_ _04091_ _04095_ _05815_ VGND VGND VPWR VPWR _02600_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15734_ _08411_ _03215_ _03223_ _02993_ VGND VGND VPWR VPWR _03224_ sky130_fd_sc_hd__a31o_1
X_12946_ _07256_ VGND VGND VPWR VPWR _07387_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_153_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15214__125 clknet_1_1__leaf__02752_ VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__inv_2
XFILLER_0_158_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15665_ _02936_ _03149_ _03156_ _02934_ VGND VGND VPWR VPWR _03157_ sky130_fd_sc_hd__o211a_1
X_12877_ CPU.registerFile\[1\]\[1\] _07255_ _07317_ _07318_ VGND VGND VPWR VPWR _07319_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_150 _07268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_161 _07322_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_172 _07412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17404_ net593 _01692_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_bitcount\[4\] sky130_fd_sc_hd__dfxtp_1
X_11828_ net2365 _05675_ _06675_ VGND VGND VPWR VPWR _06678_ sky130_fd_sc_hd__mux2_1
XANTENNA_183 _07601_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15596_ CPU.registerFile\[9\]\[6\] _02778_ _02780_ VGND VGND VPWR VPWR _03089_ sky130_fd_sc_hd__o21a_1
XANTENNA_194 _07841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17335_ net524 _01623_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11759_ _06641_ VGND VGND VPWR VPWR _01686_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17266_ net456 _01554_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload103 clknet_1_0__leaf__07223_ VGND VGND VPWR VPWR clkload103/X sky130_fd_sc_hd__clkbuf_8
X_16217_ CPU.registerFile\[28\]\[23\] CPU.registerFile\[24\]\[23\] _02772_ VGND VGND
+ VPWR VPWR _03693_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload114 clknet_1_0__leaf__03968_ VGND VGND VPWR VPWR clkload114/Y sky130_fd_sc_hd__clkinvlp_4
X_13429_ CPU.registerFile\[29\]\[15\] _07556_ _07557_ CPU.registerFile\[25\]\[15\]
+ _07856_ VGND VGND VPWR VPWR _07857_ sky130_fd_sc_hd__o221a_1
Xclkbuf_1_1__f__08431_ clknet_0__08431_ VGND VGND VPWR VPWR clknet_1_1__leaf__08431_
+ sky130_fd_sc_hd__clkbuf_16
X_17197_ clknet_leaf_11_clk _01485_ VGND VGND VPWR VPWR CPU.Bimm\[7\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_102_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__08462_ _08462_ VGND VGND VPWR VPWR clknet_0__08462_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_51_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16148_ CPU.registerFile\[22\]\[21\] CPU.registerFile\[23\]\[21\] _03066_ VGND VGND
+ VPWR VPWR _03626_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__08362_ clknet_0__08362_ VGND VGND VPWR VPWR clknet_1_1__leaf__08362_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16079_ CPU.registerFile\[28\]\[19\] CPU.registerFile\[24\]\[19\] _02761_ VGND VGND
+ VPWR VPWR _03559_ sky130_fd_sc_hd__mux2_1
X_08970_ _04688_ VGND VGND VPWR VPWR _04689_ sky130_fd_sc_hd__clkbuf_4
X_16924__4 clknet_1_1__leaf__07220_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__inv_2
XFILLER_0_127_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput1 RXD VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09522_ _04672_ _05216_ _05219_ _04679_ VGND VGND VPWR VPWR _05220_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_84_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09453_ _04716_ _05153_ _04717_ VGND VGND VPWR VPWR _05154_ sky130_fd_sc_hd__o21a_1
X_15189__102 clknet_1_0__leaf__02750_ VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__inv_2
XFILLER_0_148_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09384_ _05083_ _05073_ _05072_ _05088_ VGND VGND VPWR VPWR _05089_ sky130_fd_sc_hd__or4b_4
XFILLER_0_47_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14336__476 clknet_1_1__leaf__08466_ VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__inv_2
XFILLER_0_113_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_131_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13974__258 clknet_1_0__leaf__08357_ VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__inv_2
X_10090_ net1625 _04933_ _05633_ VGND VGND VPWR VPWR _05642_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15024__1096 clknet_1_0__leaf__02717_ VGND VGND VPWR VPWR net1128 sky130_fd_sc_hd__inv_2
X_12800_ CPU.registerFile\[23\]\[0\] _07236_ _07239_ CPU.registerFile\[19\]\[0\] _07242_
+ VGND VGND VPWR VPWR _07243_ sky130_fd_sc_hd__o221a_1
X_13780_ CPU.registerFile\[8\]\[26\] CPU.registerFile\[12\]\[26\] _05283_ VGND VGND
+ VPWR VPWR _08197_ sky130_fd_sc_hd__mux2_1
X_10992_ net2203 _05706_ _06190_ VGND VGND VPWR VPWR _06198_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14802__896 clknet_1_1__leaf__02695_ VGND VGND VPWR VPWR net928 sky130_fd_sc_hd__inv_2
XFILLER_0_69_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12731_ _07210_ VGND VGND VPWR VPWR _01258_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14046__322 clknet_1_0__leaf__08365_ VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__inv_2
X_15450_ _02936_ _02946_ VGND VGND VPWR VPWR _02947_ sky130_fd_sc_hd__or2_1
X_14501__624 clknet_1_1__leaf__02666_ VGND VGND VPWR VPWR net656 sky130_fd_sc_hd__inv_2
XFILLER_0_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12662_ CPU.cycles\[18\] _07156_ VGND VGND VPWR VPWR _07158_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11613_ net1373 _06494_ _06545_ _06539_ VGND VGND VPWR VPWR _01735_ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15381_ _02809_ VGND VGND VPWR VPWR _02879_ sky130_fd_sc_hd__buf_4
X_12593_ net1328 VGND VGND VPWR VPWR _00015_ sky130_fd_sc_hd__inv_2
X_12777__226 clknet_1_0__leaf__07225_ VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__inv_2
XFILLER_0_65_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17120_ clknet_leaf_18_clk _00022_ VGND VGND VPWR VPWR CPU.cycles\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11544_ net1393 _06495_ _06498_ _06006_ VGND VGND VPWR VPWR _01757_ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17051_ net309 _01373_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_14263_ _05054_ _05080_ _05100_ _08441_ VGND VGND VPWR VPWR _08442_ sky130_fd_sc_hd__or4_1
X_11475_ _06454_ VGND VGND VPWR VPWR _01786_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16002_ CPU.registerFile\[9\]\[17\] _08404_ _05071_ VGND VGND VPWR VPWR _03484_ sky130_fd_sc_hd__o21a_1
X_13214_ _05284_ VGND VGND VPWR VPWR _07648_ sky130_fd_sc_hd__buf_4
X_10426_ mapped_spi_flash.cmd_addr\[21\] _05825_ _05827_ mapped_spi_flash.cmd_addr\[22\]
+ VGND VGND VPWR VPWR _05847_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13145_ CPU.registerFile\[2\]\[7\] _07388_ VGND VGND VPWR VPWR _07581_ sky130_fd_sc_hd__or2_1
Xclkbuf_0__02671_ _02671_ VGND VGND VPWR VPWR clknet_0__02671_ sky130_fd_sc_hd__clkbuf_16
X_10357_ _05800_ VGND VGND VPWR VPWR _02250_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13076_ _07359_ VGND VGND VPWR VPWR _07514_ sky130_fd_sc_hd__buf_6
X_17953_ net1141 _02237_ VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dfxtp_1
X_10288_ _05763_ VGND VGND VPWR VPWR _02297_ sky130_fd_sc_hd__clkbuf_1
X_12027_ _06782_ VGND VGND VPWR VPWR _06783_ sky130_fd_sc_hd__buf_4
X_16904_ CPU.mem_wdata\[3\] _04174_ _04179_ _04176_ VGND VGND VPWR VPWR _02637_ sky130_fd_sc_hd__o211a_1
X_17884_ net1073 net1471 VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[2\] sky130_fd_sc_hd__dfxtp_1
X_16835_ per_uart.uart0.tx_bitcount\[3\] _04131_ VGND VGND VPWR VPWR _04134_ sky130_fd_sc_hd__xor2_1
XFILLER_0_73_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16766_ _04032_ net1544 VGND VGND VPWR VPWR _04081_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_66_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12929_ _05337_ VGND VGND VPWR VPWR _07370_ sky130_fd_sc_hd__clkbuf_4
X_15717_ _03200_ _03206_ _02879_ VGND VGND VPWR VPWR _03207_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_66_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16697_ _08379_ _05259_ _04006_ VGND VGND VPWR VPWR _04023_ sky130_fd_sc_hd__or3b_1
XFILLER_0_87_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14777__873 clknet_1_1__leaf__02693_ VGND VGND VPWR VPWR net905 sky130_fd_sc_hd__inv_2
X_15648_ _05406_ VGND VGND VPWR VPWR _03140_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_158_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18367_ clknet_leaf_9_clk _02645_ VGND VGND VPWR VPWR per_uart.d_in_uart\[7\] sky130_fd_sc_hd__dfxtp_1
X_15579_ CPU.registerFile\[22\]\[5\] CPU.registerFile\[23\]\[5\] _02828_ VGND VGND
+ VPWR VPWR _03073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17318_ net507 _01606_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18298_ net131 _02578_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15056__1122 clknet_1_1__leaf__02722_ VGND VGND VPWR VPWR net1154 sky130_fd_sc_hd__inv_2
X_17249_ net439 _01537_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08953_ _04671_ VGND VGND VPWR VPWR _04672_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08884_ CPU.PC\[17\] _04598_ _04602_ _04603_ VGND VGND VPWR VPWR _04604_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Left_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__02660_ clknet_0__02660_ VGND VGND VPWR VPWR clknet_1_0__leaf__02660_
+ sky130_fd_sc_hd__clkbuf_16
X_09505_ _05201_ _05203_ _04670_ VGND VGND VPWR VPWR _05204_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09436_ _04923_ _05137_ VGND VGND VPWR VPWR _05138_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09367_ _04504_ _05071_ _04777_ VGND VGND VPWR VPWR _05072_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09298_ _05000_ _04990_ _04988_ _05006_ VGND VGND VPWR VPWR _05007_ sky130_fd_sc_hd__or4b_4
XANTENNA_50 _04762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_25_Left_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_61 _05046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 _05149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_83 _05229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_94 _05332_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11260_ _06340_ VGND VGND VPWR VPWR _01887_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15243__151 clknet_1_1__leaf__02755_ VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__inv_2
X_10211_ _05229_ VGND VGND VPWR VPWR _05717_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11191_ _05520_ net1952 _06299_ VGND VGND VPWR VPWR _06304_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10142_ _05594_ _05669_ VGND VGND VPWR VPWR _05670_ sky130_fd_sc_hd__nor2_2
X_10073_ _05632_ VGND VGND VPWR VPWR _05633_ sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_34_Left_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_128_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13901_ CPU.registerFile\[13\]\[30\] _07361_ _07283_ CPU.registerFile\[9\]\[30\]
+ _07554_ VGND VGND VPWR VPWR _08314_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_145_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13832_ CPU.registerFile\[31\]\[28\] _07772_ _07773_ CPU.registerFile\[27\]\[28\]
+ _08246_ VGND VGND VPWR VPWR _08247_ sky130_fd_sc_hd__o221a_1
X_16620_ _03985_ VGND VGND VPWR VPWR _02547_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__08434_ clknet_0__08434_ VGND VGND VPWR VPWR clknet_1_0__leaf__08434_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_18_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13763_ _07639_ _08177_ _08178_ _08179_ _07570_ VGND VGND VPWR VPWR _08180_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_48_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10975_ net1652 _05689_ _06179_ VGND VGND VPWR VPWR _06189_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_48_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__08365_ clknet_0__08365_ VGND VGND VPWR VPWR clknet_1_0__leaf__08365_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_84_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12714_ per_uart.uart0.tx_count16\[1\] per_uart.uart0.tx_count16\[0\] VGND VGND VPWR
+ VPWR _07196_ sky130_fd_sc_hd__or2_1
X_15502_ CPU.registerFile\[8\]\[4\] CPU.registerFile\[12\]\[4\] _02852_ VGND VGND
+ VPWR VPWR _02997_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16482_ _02924_ _03947_ _03948_ _03949_ _02782_ VGND VGND VPWR VPWR _03950_ sky130_fd_sc_hd__a221o_1
XFILLER_0_155_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13694_ CPU.registerFile\[2\]\[24\] _07322_ VGND VGND VPWR VPWR _08113_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15433_ _05093_ VGND VGND VPWR VPWR _02930_ sky130_fd_sc_hd__buf_4
X_18221_ net62 _02501_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_12645_ CPU.cycles\[10\] CPU.cycles\[11\] _07146_ VGND VGND VPWR VPWR _07148_ sky130_fd_sc_hd__and3_1
XFILLER_0_53_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_61_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18152_ clknet_leaf_19_clk _02432_ VGND VGND VPWR VPWR CPU.aluIn1\[18\] sky130_fd_sc_hd__dfxtp_2
X_15364_ CPU.registerFile\[8\]\[1\] _02861_ VGND VGND VPWR VPWR _02862_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12576_ _07111_ VGND VGND VPWR VPWR _01271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17103_ _00013_ _00014_ VGND VGND VPWR VPWR CPU.writeBack sky130_fd_sc_hd__dlxtn_2
XFILLER_0_136_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18083_ net146 _02363_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_11527_ _06488_ VGND VGND VPWR VPWR _06489_ sky130_fd_sc_hd__buf_2
X_15295_ _08396_ VGND VGND VPWR VPWR _02794_ sky130_fd_sc_hd__buf_4
XFILLER_0_81_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17034_ net292 _01356_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[28\] sky130_fd_sc_hd__dfxtp_1
Xhold309 CPU.registerFile\[5\]\[30\] VGND VGND VPWR VPWR net1550 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11458_ _05514_ net1946 _06444_ VGND VGND VPWR VPWR _06446_ sky130_fd_sc_hd__mux2_1
X_14319__460 clknet_1_1__leaf__08465_ VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__inv_2
XFILLER_0_33_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__02723_ _02723_ VGND VGND VPWR VPWR clknet_0__02723_ sky130_fd_sc_hd__clkbuf_16
X_10409_ _05830_ _05835_ VGND VGND VPWR VPWR _05836_ sky130_fd_sc_hd__and2_1
X_14177_ _04619_ VGND VGND VPWR VPWR _08426_ sky130_fd_sc_hd__inv_2
X_11389_ _06409_ VGND VGND VPWR VPWR _01827_ sky130_fd_sc_hd__clkbuf_1
X_13957__242 clknet_1_0__leaf__08356_ VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__inv_2
Xclkbuf_0__02654_ _02654_ VGND VGND VPWR VPWR clknet_0__02654_ sky130_fd_sc_hd__clkbuf_16
X_13128_ _07271_ _07550_ _07553_ _07564_ _07306_ VGND VGND VPWR VPWR _07565_ sky130_fd_sc_hd__o311a_1
X_13059_ CPU.mem_wdata\[4\] _07358_ _07473_ _07497_ _05844_ VGND VGND VPWR VPWR _01299_
+ sky130_fd_sc_hd__o221a_1
X_17936_ net1125 _02220_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[16\] sky130_fd_sc_hd__dfxtp_1
Xhold1009 CPU.registerFile\[10\]\[16\] VGND VGND VPWR VPWR net2250 sky130_fd_sc_hd__dlygate4sd3_1
X_14018__298 clknet_1_0__leaf__08361_ VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__inv_2
X_17867_ net1056 _02151_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14211__388 clknet_1_1__leaf__08430_ VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__inv_2
X_16818_ _07178_ _07195_ _04121_ per_uart.uart0.tx_count16\[2\] VGND VGND VPWR VPWR
+ _04122_ sky130_fd_sc_hd__a22oi_1
X_17798_ net987 _02082_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_37_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16749_ _08436_ _08459_ _05095_ VGND VGND VPWR VPWR _04067_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09221_ _04932_ VGND VGND VPWR VPWR _04933_ sky130_fd_sc_hd__buf_2
XFILLER_0_44_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09152_ _04862_ _04863_ VGND VGND VPWR VPWR _04864_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15023__1095 clknet_1_0__leaf__02717_ VGND VGND VPWR VPWR net1127 sky130_fd_sc_hd__inv_2
XFILLER_0_127_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09083_ CPU.Iimm\[4\] _04498_ _04795_ _04492_ VGND VGND VPWR VPWR _04796_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold810 CPU.registerFile\[24\]\[6\] VGND VGND VPWR VPWR net2051 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold821 CPU.registerFile\[21\]\[26\] VGND VGND VPWR VPWR net2062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold832 CPU.registerFile\[21\]\[11\] VGND VGND VPWR VPWR net2073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold843 CPU.registerFile\[31\]\[14\] VGND VGND VPWR VPWR net2084 sky130_fd_sc_hd__dlygate4sd3_1
Xhold854 mapped_spi_flash.rcv_data\[19\] VGND VGND VPWR VPWR net2095 sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 CPU.registerFile\[16\]\[8\] VGND VGND VPWR VPWR net2106 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14530__650 clknet_1_1__leaf__02669_ VGND VGND VPWR VPWR net682 sky130_fd_sc_hd__inv_2
Xhold876 CPU.registerFile\[17\]\[12\] VGND VGND VPWR VPWR net2117 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__08428_ _08428_ VGND VGND VPWR VPWR clknet_0__08428_ sky130_fd_sc_hd__clkbuf_16
Xhold887 CPU.registerFile\[19\]\[31\] VGND VGND VPWR VPWR net2128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold898 CPU.registerFile\[2\]\[1\] VGND VGND VPWR VPWR net2139 sky130_fd_sc_hd__dlygate4sd3_1
X_09985_ _05585_ VGND VGND VPWR VPWR _02454_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08936_ _04504_ _04619_ _04655_ VGND VGND VPWR VPWR _04656_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_0__08359_ _08359_ VGND VGND VPWR VPWR clknet_0__08359_ sky130_fd_sc_hd__clkbuf_16
X_08867_ CPU.PC\[21\] _04586_ VGND VGND VPWR VPWR _04587_ sky130_fd_sc_hd__nand2_1
X_14448__577 clknet_1_0__leaf__02660_ VGND VGND VPWR VPWR net609 sky130_fd_sc_hd__inv_2
XFILLER_0_99_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08798_ CPU.aluIn1\[4\] net1276 VGND VGND VPWR VPWR _04518_ sky130_fd_sc_hd__nand2_1
Xclkbuf_1_0__f__02712_ clknet_0__02712_ VGND VGND VPWR VPWR clknet_1_0__leaf__02712_
+ sky130_fd_sc_hd__clkbuf_16
X_14186__365 clknet_1_0__leaf__08428_ VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__inv_2
XFILLER_0_79_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10760_ _05499_ net1749 _06070_ VGND VGND VPWR VPWR _06075_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09419_ _04437_ _04806_ _05121_ _04768_ VGND VGND VPWR VPWR _05122_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_94_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10691_ _06038_ VGND VGND VPWR VPWR _02154_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12430_ _05170_ net1973 _07024_ VGND VGND VPWR VPWR _07034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12361_ _06997_ VGND VGND VPWR VPWR _01405_ sky130_fd_sc_hd__clkbuf_1
X_14914__997 clknet_1_0__leaf__02706_ VGND VGND VPWR VPWR net1029 sky130_fd_sc_hd__inv_2
XFILLER_0_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14100_ CPU.instr\[2\] _05386_ _00000_ VGND VGND VPWR VPWR _08378_ sky130_fd_sc_hd__mux2_1
X_11312_ _05505_ net1999 _06360_ VGND VGND VPWR VPWR _06368_ sky130_fd_sc_hd__mux2_1
X_14613__725 clknet_1_0__leaf__02677_ VGND VGND VPWR VPWR net757 sky130_fd_sc_hd__inv_2
X_15080_ _04192_ _07195_ VGND VGND VPWR VPWR _02726_ sky130_fd_sc_hd__nand2_1
X_12292_ _06954_ VGND VGND VPWR VPWR _01431_ sky130_fd_sc_hd__clkbuf_1
X_14031_ clknet_1_1__leaf__07222_ VGND VGND VPWR VPWR _08363_ sky130_fd_sc_hd__buf_1
X_11243_ _06331_ VGND VGND VPWR VPWR _01895_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11174_ _05503_ net2526 _06288_ VGND VGND VPWR VPWR _06295_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_42_Left_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10125_ _05660_ VGND VGND VPWR VPWR _02357_ sky130_fd_sc_hd__clkbuf_1
X_15982_ CPU.registerFile\[5\]\[17\] CPU.registerFile\[4\]\[17\] _02898_ VGND VGND
+ VPWR VPWR _03464_ sky130_fd_sc_hd__mux2_1
X_17721_ net910 _02005_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_10056_ _05623_ VGND VGND VPWR VPWR _02389_ sky130_fd_sc_hd__clkbuf_1
X_17652_ net841 _01940_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_15055__1121 clknet_1_1__leaf__02722_ VGND VGND VPWR VPWR net1153 sky130_fd_sc_hd__inv_2
X_16603_ _03972_ _03973_ VGND VGND VPWR VPWR _03974_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13815_ _07330_ _08230_ VGND VGND VPWR VPWR _08231_ sky130_fd_sc_hd__or2_1
X_14795_ clknet_1_1__leaf__02686_ VGND VGND VPWR VPWR _02695_ sky130_fd_sc_hd__buf_1
X_17583_ net772 _01871_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13746_ _07418_ _08162_ _08163_ VGND VGND VPWR VPWR _08164_ sky130_fd_sc_hd__o21a_1
X_10958_ _06180_ VGND VGND VPWR VPWR _02029_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_51_Left_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_158_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_158_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13677_ CPU.registerFile\[3\]\[23\] _07577_ VGND VGND VPWR VPWR _08097_ sky130_fd_sc_hd__or2_1
X_16465_ _03929_ _03932_ _02858_ VGND VGND VPWR VPWR _03933_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10889_ net1700 _05668_ _06143_ VGND VGND VPWR VPWR _06144_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_158_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18204_ net45 _02484_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_15416_ CPU.registerFile\[11\]\[2\] _02895_ _02911_ _02912_ VGND VGND VPWR VPWR _02913_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12628_ net1467 _07136_ VGND VGND VPWR VPWR _07139_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16396_ CPU.registerFile\[7\]\[29\] _02898_ _02999_ _03865_ VGND VGND VPWR VPWR _03866_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_143_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15347_ _07308_ VGND VGND VPWR VPWR _02846_ sky130_fd_sc_hd__buf_2
X_18135_ clknet_leaf_28_clk _02415_ VGND VGND VPWR VPWR CPU.aluIn1\[1\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_143_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12559_ _07102_ VGND VGND VPWR VPWR _01279_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14889__974 clknet_1_0__leaf__02704_ VGND VGND VPWR VPWR net1006 sky130_fd_sc_hd__inv_2
X_18066_ net1239 _02346_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15278_ _05405_ VGND VGND VPWR VPWR _02777_ sky130_fd_sc_hd__buf_4
XFILLER_0_112_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold106 mapped_spi_flash.cmd_addr\[24\] VGND VGND VPWR VPWR net1347 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold117 mapped_spi_ram.cmd_addr\[17\] VGND VGND VPWR VPWR net1358 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold128 mapped_spi_flash.cmd_addr\[23\] VGND VGND VPWR VPWR net1369 sky130_fd_sc_hd__dlygate4sd3_1
X_17017_ net275 _01339_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold139 _07161_ VGND VGND VPWR VPWR net1380 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_655 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__02706_ _02706_ VGND VGND VPWR VPWR clknet_0__02706_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_107_Right_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09770_ _05455_ VGND VGND VPWR VPWR _02539_ sky130_fd_sc_hd__clkbuf_1
X_08721_ _04392_ _04440_ _04333_ VGND VGND VPWR VPWR _04441_ sky130_fd_sc_hd__o21a_1
X_17919_ net1108 _02203_ VGND VGND VPWR VPWR mapped_spi_flash.snd_bitcount\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08652_ CPU.instr\[5\] VGND VGND VPWR VPWR _04372_ sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_1_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08583_ _04297_ _04299_ _04290_ VGND VGND VPWR VPWR _04303_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_105_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09204_ _04915_ VGND VGND VPWR VPWR _04916_ sky130_fd_sc_hd__buf_2
XFILLER_0_119_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09135_ CPU.Jimm\[13\] _04829_ _04831_ VGND VGND VPWR VPWR _04847_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09066_ _04779_ VGND VGND VPWR VPWR _04780_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold640 CPU.registerFile\[2\]\[28\] VGND VGND VPWR VPWR net1881 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold651 CPU.registerFile\[14\]\[3\] VGND VGND VPWR VPWR net1892 sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 CPU.registerFile\[14\]\[8\] VGND VGND VPWR VPWR net1903 sky130_fd_sc_hd__dlygate4sd3_1
Xhold673 CPU.registerFile\[13\]\[17\] VGND VGND VPWR VPWR net1914 sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 CPU.registerFile\[3\]\[25\] VGND VGND VPWR VPWR net1925 sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 CPU.registerFile\[2\]\[20\] VGND VGND VPWR VPWR net1936 sky130_fd_sc_hd__dlygate4sd3_1
X_09968_ _05576_ VGND VGND VPWR VPWR _02462_ sky130_fd_sc_hd__clkbuf_1
X_08919_ CPU.PC\[2\] _04598_ _04638_ _04626_ VGND VGND VPWR VPWR _04639_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_125_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09899_ _05534_ VGND VGND VPWR VPWR _02489_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_525 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11930_ _06731_ VGND VGND VPWR VPWR _01605_ sky130_fd_sc_hd__clkbuf_1
X_11861_ net2352 _05708_ _06686_ VGND VGND VPWR VPWR _06695_ sky130_fd_sc_hd__mux2_1
X_13600_ CPU.registerFile\[14\]\[21\] CPU.registerFile\[10\]\[21\] _04936_ VGND VGND
+ VPWR VPWR _08022_ sky130_fd_sc_hd__mux2_1
X_10812_ _05551_ net1697 _06092_ VGND VGND VPWR VPWR _06102_ sky130_fd_sc_hd__mux2_1
X_11792_ _06658_ VGND VGND VPWR VPWR _01670_ sky130_fd_sc_hd__clkbuf_1
X_13531_ _07364_ _07954_ VGND VGND VPWR VPWR _07955_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_844 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10743_ _06065_ VGND VGND VPWR VPWR _02129_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16250_ CPU.registerFile\[22\]\[24\] CPU.registerFile\[23\]\[24\] _03066_ VGND VGND
+ VPWR VPWR _03725_ sky130_fd_sc_hd__mux2_1
X_13462_ CPU.registerFile\[14\]\[16\] CPU.registerFile\[10\]\[16\] _07492_ VGND VGND
+ VPWR VPWR _07889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10674_ mapped_spi_flash.rcv_bitcount\[1\] mapped_spi_flash.rcv_bitcount\[0\] VGND
+ VGND VPWR VPWR _06028_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12413_ _07025_ VGND VGND VPWR VPWR _01381_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16181_ CPU.registerFile\[7\]\[22\] _03317_ VGND VGND VPWR VPWR _03658_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13393_ _07818_ _07819_ _07821_ VGND VGND VPWR VPWR _07822_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_153_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12344_ _04982_ net1789 _06988_ VGND VGND VPWR VPWR _06989_ sky130_fd_sc_hd__mux2_1
X_12275_ CPU.aluReg\[11\] _06941_ _06924_ VGND VGND VPWR VPWR _06942_ sky130_fd_sc_hd__mux2_1
X_11226_ _05555_ net1873 _06287_ VGND VGND VPWR VPWR _06322_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11157_ _06285_ VGND VGND VPWR VPWR _01935_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10108_ _05651_ VGND VGND VPWR VPWR _02365_ sky130_fd_sc_hd__clkbuf_1
X_11088_ _06248_ VGND VGND VPWR VPWR _01967_ sky130_fd_sc_hd__clkbuf_1
X_15965_ _03443_ _03447_ _03138_ VGND VGND VPWR VPWR _03448_ sky130_fd_sc_hd__a21o_1
X_17704_ net893 _01992_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_10039_ _05614_ VGND VGND VPWR VPWR _02397_ sky130_fd_sc_hd__clkbuf_1
X_15022__1094 clknet_1_0__leaf__02717_ VGND VGND VPWR VPWR net1126 sky130_fd_sc_hd__inv_2
X_15896_ CPU.registerFile\[25\]\[14\] _03280_ _02803_ VGND VGND VPWR VPWR _03381_
+ sky130_fd_sc_hd__o21a_1
X_17635_ net824 _01923_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_17566_ net755 _01854_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13729_ CPU.registerFile\[17\]\[25\] _07480_ _07305_ VGND VGND VPWR VPWR _08147_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17497_ net686 _01785_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16448_ CPU.registerFile\[27\]\[30\] _02889_ _02780_ VGND VGND VPWR VPWR _03917_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16379_ CPU.registerFile\[6\]\[28\] CPU.registerFile\[7\]\[28\] _02819_ VGND VGND
+ VPWR VPWR _03850_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18118_ net181 _02398_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18049_ net1222 _02329_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09822_ _05482_ VGND VGND VPWR VPWR _02514_ sky130_fd_sc_hd__clkbuf_1
X_09753_ _05232_ _05235_ _04636_ VGND VGND VPWR VPWR _05442_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08704_ _04313_ _04273_ VGND VGND VPWR VPWR _04424_ sky130_fd_sc_hd__or2b_1
X_09684_ _04871_ _04876_ _04877_ VGND VGND VPWR VPWR _05376_ sky130_fd_sc_hd__nand3_1
XFILLER_0_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14642__751 clknet_1_0__leaf__02680_ VGND VGND VPWR VPWR net783 sky130_fd_sc_hd__inv_2
X_08635_ CPU.aluIn1\[26\] _04231_ VGND VGND VPWR VPWR _04355_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_87_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ CPU.mem_wdata\[3\] CPU.Iimm\[3\] _04202_ VGND VGND VPWR VPWR _04286_ sky130_fd_sc_hd__mux2_2
XFILLER_0_77_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08497_ _04216_ _04208_ VGND VGND VPWR VPWR _04217_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14040__317 clknet_1_0__leaf__08364_ VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__inv_2
XFILLER_0_44_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09118_ CPU.instr\[3\] _04292_ VGND VGND VPWR VPWR _04830_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_118_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10390_ _05817_ VGND VGND VPWR VPWR _05820_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_135_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15054__1120 clknet_1_1__leaf__02722_ VGND VGND VPWR VPWR net1152 sky130_fd_sc_hd__inv_2
X_09049_ _04763_ VGND VGND VPWR VPWR _02576_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12060_ _06800_ VGND VGND VPWR VPWR _01543_ sky130_fd_sc_hd__clkbuf_1
Xhold470 CPU.registerFile\[5\]\[27\] VGND VGND VPWR VPWR net1711 sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 CPU.registerFile\[30\]\[0\] VGND VGND VPWR VPWR net1722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold492 CPU.registerFile\[12\]\[21\] VGND VGND VPWR VPWR net1733 sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ net2311 _05725_ _06201_ VGND VGND VPWR VPWR _06208_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_8_Left_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14725__826 clknet_1_1__leaf__02688_ VGND VGND VPWR VPWR net858 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_51_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12962_ _07402_ VGND VGND VPWR VPWR _07403_ sky130_fd_sc_hd__clkbuf_8
X_15750_ _02901_ _03237_ _03238_ _02867_ VGND VGND VPWR VPWR _03239_ sky130_fd_sc_hd__a22o_1
Xhold1170 CPU.registerFile\[8\]\[15\] VGND VGND VPWR VPWR net2411 sky130_fd_sc_hd__dlygate4sd3_1
X_11913_ net2536 _05691_ _06722_ VGND VGND VPWR VPWR _06723_ sky130_fd_sc_hd__mux2_1
Xhold1181 CPU.registerFile\[2\]\[6\] VGND VGND VPWR VPWR net2422 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1192 CPU.aluIn1\[27\] VGND VGND VPWR VPWR net2433 sky130_fd_sc_hd__dlygate4sd3_1
X_12893_ _07321_ _07333_ _07334_ VGND VGND VPWR VPWR _07335_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15681_ CPU.registerFile\[27\]\[8\] CPU.registerFile\[31\]\[8\] _03050_ VGND VGND
+ VPWR VPWR _03172_ sky130_fd_sc_hd__mux2_1
XANTENNA_310 _07914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_321 _07914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17420_ net609 _01708_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[13\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_332 CPU.mem_wdata\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11844_ _06674_ VGND VGND VPWR VPWR _06686_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_343 _05071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_354 _07268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_365 _02889_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_376 _07291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17351_ net540 _01639_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[15\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_387 _07250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11775_ _06649_ VGND VGND VPWR VPWR _01678_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_398 _07250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_155_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ CPU.registerFile\[2\]\[26\] _02872_ _02873_ CPU.registerFile\[3\]\[26\] _02875_
+ VGND VGND VPWR VPWR _03775_ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13514_ CPU.registerFile\[14\]\[18\] CPU.registerFile\[10\]\[18\] _07476_ VGND VGND
+ VPWR VPWR _07939_ sky130_fd_sc_hd__mux2_1
X_10726_ _05532_ net1578 _06056_ VGND VGND VPWR VPWR _06057_ sky130_fd_sc_hd__mux2_1
X_17282_ net471 _01570_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13445_ CPU.registerFile\[1\]\[16\] _07576_ _07871_ _07639_ VGND VGND VPWR VPWR _07872_
+ sky130_fd_sc_hd__a22o_1
X_16233_ CPU.registerFile\[28\]\[24\] _03064_ VGND VGND VPWR VPWR _03708_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14771__868 clknet_1_1__leaf__02692_ VGND VGND VPWR VPWR net900 sky130_fd_sc_hd__inv_2
XFILLER_0_152_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10657_ mapped_spi_flash.state\[0\] mapped_spi_flash.state\[3\] VGND VGND VPWR VPWR
+ _06015_ sky130_fd_sc_hd__nor2_1
Xclkload15 clknet_leaf_18_clk VGND VGND VPWR VPWR clkload15/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload26 clknet_leaf_10_clk VGND VGND VPWR VPWR clkload26/Y sky130_fd_sc_hd__clkinv_4
X_16531__198 clknet_1_0__leaf__03964_ VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__inv_2
XFILLER_0_106_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13376_ CPU.registerFile\[3\]\[14\] _07804_ _07376_ VGND VGND VPWR VPWR _07805_ sky130_fd_sc_hd__o21a_1
XFILLER_0_24_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload37 clknet_1_0__leaf__02720_ VGND VGND VPWR VPWR clkload37/X sky130_fd_sc_hd__clkbuf_8
X_16164_ CPU.registerFile\[30\]\[22\] CPU.registerFile\[26\]\[22\] _02918_ VGND VGND
+ VPWR VPWR _03641_ sky130_fd_sc_hd__mux2_1
X_10588_ net1468 _05968_ _05975_ _05936_ VGND VGND VPWR VPWR _02193_ sky130_fd_sc_hd__o211a_1
Xclkload48 clknet_1_1__leaf__02716_ VGND VGND VPWR VPWR clkload48/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload59 clknet_1_1__leaf__02696_ VGND VGND VPWR VPWR clkload59/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_106_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12327_ _04714_ net2067 _06977_ VGND VGND VPWR VPWR _06980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16095_ _03022_ _03571_ _03572_ _03573_ _03028_ VGND VGND VPWR VPWR _03574_ sky130_fd_sc_hd__o221a_1
X_12258_ CPU.aluReg\[15\] _06928_ _06924_ VGND VGND VPWR VPWR _06929_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11209_ _06313_ VGND VGND VPWR VPWR _01911_ sky130_fd_sc_hd__clkbuf_1
X_12189_ net2452 _06875_ _06862_ VGND VGND VPWR VPWR _06876_ sky130_fd_sc_hd__mux2_1
X_16997_ clknet_leaf_21_clk _01323_ VGND VGND VPWR VPWR CPU.rs2\[28\] sky130_fd_sc_hd__dfxtp_1
X_14364__501 clknet_1_0__leaf__02652_ VGND VGND VPWR VPWR net533 sky130_fd_sc_hd__inv_2
X_15948_ CPU.registerFile\[14\]\[16\] CPU.registerFile\[10\]\[16\] _03082_ VGND VGND
+ VPWR VPWR _03431_ sky130_fd_sc_hd__mux2_1
X_15879_ _02757_ _03341_ _03350_ _03364_ _02846_ VGND VGND VPWR VPWR _03365_ sky130_fd_sc_hd__a311o_2
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_69_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17618_ net807 _01906_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_102_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17549_ net738 _01837_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload9 clknet_leaf_12_clk VGND VGND VPWR VPWR clkload9/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_132_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09805_ _05473_ VGND VGND VPWR VPWR _02522_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09736_ _05425_ VGND VGND VPWR VPWR _05426_ sky130_fd_sc_hd__clkbuf_4
X_09667_ net1638 _05359_ _05189_ VGND VGND VPWR VPWR _05360_ sky130_fd_sc_hd__mux2_1
X_08618_ _04337_ VGND VGND VPWR VPWR _04338_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09598_ _04864_ _04882_ VGND VGND VPWR VPWR _05293_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08549_ CPU.aluIn1\[9\] _04268_ VGND VGND VPWR VPWR _04269_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11560_ _06501_ _05882_ VGND VGND VPWR VPWR _06510_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10511_ _04516_ _05914_ _05916_ VGND VGND VPWR VPWR _05917_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11491_ _05547_ net1917 _06455_ VGND VGND VPWR VPWR _06463_ sky130_fd_sc_hd__mux2_1
X_13230_ _07418_ _07662_ _07663_ VGND VGND VPWR VPWR _07664_ sky130_fd_sc_hd__o21a_1
X_10442_ net1401 _05850_ _05851_ _05859_ VGND VGND VPWR VPWR _05860_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_133_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15021__1093 clknet_1_0__leaf__02717_ VGND VGND VPWR VPWR net1125 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_150_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13161_ CPU.registerFile\[14\]\[7\] CPU.registerFile\[10\]\[7\] _07492_ VGND VGND
+ VPWR VPWR _07597_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10373_ _05808_ VGND VGND VPWR VPWR _02242_ sky130_fd_sc_hd__clkbuf_1
X_12112_ _04933_ net2145 _06819_ VGND VGND VPWR VPWR _06828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13092_ _07525_ _07526_ _07527_ _07529_ _07302_ VGND VGND VPWR VPWR _07530_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_53_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12043_ _06791_ VGND VGND VPWR VPWR _01551_ sky130_fd_sc_hd__clkbuf_1
X_16920_ net2262 _04182_ VGND VGND VPWR VPWR _04189_ sky130_fd_sc_hd__or2_1
X_14313__455 clknet_1_0__leaf__08464_ VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__inv_2
X_16851_ net1565 per_uart.rx_data\[4\] _04139_ VGND VGND VPWR VPWR _04144_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_148_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13951__237 clknet_1_0__leaf__07226_ VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__inv_2
X_15802_ CPU.registerFile\[20\]\[11\] CPU.registerFile\[21\]\[11\] _03066_ VGND VGND
+ VPWR VPWR _03290_ sky130_fd_sc_hd__mux2_1
X_16782_ _04050_ _04092_ _04093_ _04094_ VGND VGND VPWR VPWR _04095_ sky130_fd_sc_hd__a31o_1
X_15733_ _02903_ _03219_ _03222_ VGND VGND VPWR VPWR _03223_ sky130_fd_sc_hd__or3_1
X_12945_ CPU.registerFile\[21\]\[2\] _07382_ _07383_ CPU.registerFile\[17\]\[2\] _07385_
+ VGND VGND VPWR VPWR _07386_ sky130_fd_sc_hd__o221a_1
XFILLER_0_62_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15664_ _02948_ _03152_ _03155_ VGND VGND VPWR VPWR _03156_ sky130_fd_sc_hd__or3_2
XANTENNA_140 _05702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12876_ _05284_ VGND VGND VPWR VPWR _07318_ sky130_fd_sc_hd__buf_6
XANTENNA_151 _07268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_162 _07322_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17403_ net592 _01691_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_bitcount\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_173 _07433_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11827_ _06677_ VGND VGND VPWR VPWR _01654_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_184 _07621_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15595_ CPU.registerFile\[13\]\[6\] _02775_ VGND VGND VPWR VPWR _03088_ sky130_fd_sc_hd__or2_1
XANTENNA_195 _07841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17334_ net523 _01622_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_11758_ _04696_ net1915 _06639_ VGND VGND VPWR VPWR _06641_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_778 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10709_ _05516_ net2417 _06045_ VGND VGND VPWR VPWR _06048_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17265_ net455 _01553_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_11689_ net1534 _06590_ _06597_ _06594_ VGND VGND VPWR VPWR _01711_ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload104 clknet_1_0__leaf__08362_ VGND VGND VPWR VPWR clkload104/Y sky130_fd_sc_hd__clkinvlp_4
X_16216_ CPU.registerFile\[30\]\[23\] CPU.registerFile\[26\]\[23\] _03247_ VGND VGND
+ VPWR VPWR _03692_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__08430_ clknet_0__08430_ VGND VGND VPWR VPWR clknet_1_1__leaf__08430_
+ sky130_fd_sc_hd__clkbuf_16
Xclkload115 clknet_1_1__leaf__03967_ VGND VGND VPWR VPWR clkload115/Y sky130_fd_sc_hd__clkinvlp_4
X_13428_ _07291_ _07855_ VGND VGND VPWR VPWR _07856_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17196_ clknet_leaf_11_clk _01484_ VGND VGND VPWR VPWR CPU.Bimm\[6\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_102_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__08361_ clknet_0__08361_ VGND VGND VPWR VPWR clknet_1_1__leaf__08361_
+ sky130_fd_sc_hd__clkbuf_16
X_13359_ CPU.registerFile\[16\]\[13\] CPU.registerFile\[20\]\[13\] _07318_ VGND VGND
+ VPWR VPWR _07789_ sky130_fd_sc_hd__mux2_1
X_16147_ _03065_ _03623_ _03624_ VGND VGND VPWR VPWR _03625_ sky130_fd_sc_hd__o21a_1
XFILLER_0_141_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16078_ _03015_ _03555_ _03556_ _03557_ _02930_ VGND VGND VPWR VPWR _03558_ sky130_fd_sc_hd__a221o_1
XFILLER_0_121_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14708__810 clknet_1_0__leaf__02687_ VGND VGND VPWR VPWR net842 sky130_fd_sc_hd__inv_2
X_14288__432 clknet_1_1__leaf__08462_ VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__inv_2
Xinput2 resetn VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_4
XFILLER_0_127_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09521_ _04672_ _05218_ VGND VGND VPWR VPWR _05219_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_84_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09452_ _04718_ _05152_ _05112_ VGND VGND VPWR VPWR _05153_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09383_ _04818_ _05085_ _05087_ _04916_ VGND VGND VPWR VPWR _05088_ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14754__852 clknet_1_0__leaf__02691_ VGND VGND VPWR VPWR net884 sky130_fd_sc_hd__inv_2
XFILLER_0_47_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16514__182 clknet_1_1__leaf__03963_ VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__inv_2
XFILLER_0_7_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_115_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_89_Left_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_98_Left_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09719_ _05406_ _05281_ _05408_ _05286_ VGND VGND VPWR VPWR _05409_ sky130_fd_sc_hd__o211a_1
X_10991_ _06197_ VGND VGND VPWR VPWR _02013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12730_ _07209_ net1597 _07205_ VGND VGND VPWR VPWR _07210_ sky130_fd_sc_hd__mux2_1
X_14837__927 clknet_1_1__leaf__02699_ VGND VGND VPWR VPWR net959 sky130_fd_sc_hd__inv_2
X_12661_ _07156_ net1417 VGND VGND VPWR VPWR _00023_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11612_ net1387 _06501_ _06496_ CPU.mem_wdata\[2\] _06508_ VGND VGND VPWR VPWR _06545_
+ sky130_fd_sc_hd__a221o_1
X_12592_ _07119_ VGND VGND VPWR VPWR _01263_ sky130_fd_sc_hd__clkbuf_1
X_15380_ _08401_ _02869_ _02877_ _02844_ VGND VGND VPWR VPWR _02878_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_873 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11543_ _06496_ _06497_ _06494_ VGND VGND VPWR VPWR _06498_ sky130_fd_sc_hd__o21ai_1
X_14262_ _05120_ _05145_ _05161_ _08440_ VGND VGND VPWR VPWR _08441_ sky130_fd_sc_hd__or4_1
X_17050_ net308 _01372_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_11474_ _05530_ net2423 _06444_ VGND VGND VPWR VPWR _06454_ sky130_fd_sc_hd__mux2_1
X_13213_ _07254_ _07640_ _07645_ _07646_ VGND VGND VPWR VPWR _07647_ sky130_fd_sc_hd__o211a_1
X_16001_ CPU.registerFile\[15\]\[17\] CPU.registerFile\[11\]\[17\] _03247_ VGND VGND
+ VPWR VPWR _03483_ sky130_fd_sc_hd__mux2_1
X_10425_ _05846_ VGND VGND VPWR VPWR _02227_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13144_ CPU.registerFile\[6\]\[7\] CPU.registerFile\[7\]\[7\] _07371_ VGND VGND VPWR
+ VPWR _07580_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__02670_ _02670_ VGND VGND VPWR VPWR clknet_0__02670_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_103_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10356_ _05532_ net2073 _05799_ VGND VGND VPWR VPWR _05800_ sky130_fd_sc_hd__mux2_1
XFILLER_0_148_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14883__969 clknet_1_1__leaf__02703_ VGND VGND VPWR VPWR net1001 sky130_fd_sc_hd__inv_2
XFILLER_0_130_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13075_ _07510_ _07512_ _07320_ VGND VGND VPWR VPWR _07513_ sky130_fd_sc_hd__mux2_1
X_17952_ clknet_leaf_22_clk _02236_ VGND VGND VPWR VPWR CPU.aluWr sky130_fd_sc_hd__dfxtp_1
X_15220__130 clknet_1_1__leaf__02753_ VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__inv_2
X_10287_ _05532_ net2188 _05762_ VGND VGND VPWR VPWR _05763_ sky130_fd_sc_hd__mux2_1
X_12026_ _05557_ _06395_ VGND VGND VPWR VPWR _06782_ sky130_fd_sc_hd__nand2_2
X_16903_ net2222 _04177_ VGND VGND VPWR VPWR _04179_ sky130_fd_sc_hd__or2_1
X_17883_ net1072 _02167_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[1\] sky130_fd_sc_hd__dfxtp_1
X_17481__27 VGND VGND VPWR VPWR _17481__27/HI net27 sky130_fd_sc_hd__conb_1
X_16834_ _05816_ net20 _04133_ _04126_ net2340 VGND VGND VPWR VPWR _02613_ sky130_fd_sc_hd__a32o_1
XFILLER_0_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_26 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16765_ _04076_ _04080_ _05942_ VGND VGND VPWR VPWR _02597_ sky130_fd_sc_hd__o21a_1
XFILLER_0_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15716_ _08401_ _03202_ _03205_ _02844_ VGND VGND VPWR VPWR _03206_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_66_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12928_ _07368_ VGND VGND VPWR VPWR _07369_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_66_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16696_ _08436_ _08459_ _05257_ VGND VGND VPWR VPWR _04022_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15647_ _03133_ _03137_ _03138_ VGND VGND VPWR VPWR _03139_ sky130_fd_sc_hd__a21o_1
X_12859_ _04785_ VGND VGND VPWR VPWR _07302_ sky130_fd_sc_hd__buf_4
XFILLER_0_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14476__602 clknet_1_1__leaf__02663_ VGND VGND VPWR VPWR net634 sky130_fd_sc_hd__inv_2
XFILLER_0_139_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18366_ clknet_leaf_9_clk _02644_ VGND VGND VPWR VPWR per_uart.d_in_uart\[6\] sky130_fd_sc_hd__dfxtp_1
X_15578_ _02791_ VGND VGND VPWR VPWR _03072_ sky130_fd_sc_hd__buf_4
XFILLER_0_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17317_ net506 _01605_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14529_ clknet_1_0__leaf__02664_ VGND VGND VPWR VPWR _02669_ sky130_fd_sc_hd__buf_1
X_18297_ net130 _02577_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17248_ net438 _01536_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_910 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17179_ clknet_leaf_12_clk _01467_ VGND VGND VPWR VPWR CPU.Bimm\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08952_ _04670_ VGND VGND VPWR VPWR _04671_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_110_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__02699_ clknet_0__02699_ VGND VGND VPWR VPWR clknet_1_1__leaf__02699_
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f__07226_ clknet_0__07226_ VGND VGND VPWR VPWR clknet_1_1__leaf__07226_
+ sky130_fd_sc_hd__clkbuf_16
X_08883_ _04559_ _04562_ _04563_ _04506_ VGND VGND VPWR VPWR _04603_ sky130_fd_sc_hd__a31o_1
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15020__1092 clknet_1_1__leaf__02717_ VGND VGND VPWR VPWR net1124 sky130_fd_sc_hd__inv_2
XFILLER_0_79_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09504_ _04267_ _05202_ VGND VGND VPWR VPWR _05203_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09435_ CPU.PC\[12\] _04922_ CPU.PC\[13\] VGND VGND VPWR VPWR _05137_ sky130_fd_sc_hd__a21oi_1
X_09366_ _05070_ VGND VGND VPWR VPWR _05071_ sky130_fd_sc_hd__buf_4
X_14342__481 clknet_1_0__leaf__08467_ VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__inv_2
XFILLER_0_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_40 _03564_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09297_ _04818_ _05003_ _05005_ _04955_ VGND VGND VPWR VPWR _05006_ sky130_fd_sc_hd__o22a_1
XFILLER_0_35_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13980__263 clknet_1_1__leaf__08358_ VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__inv_2
XFILLER_0_117_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_51 _04762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_62 _05046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_73 _05149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_84 _05229_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_95 _05332_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10210_ _05716_ VGND VGND VPWR VPWR _02328_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11190_ _06303_ VGND VGND VPWR VPWR _01920_ sky130_fd_sc_hd__clkbuf_1
X_10141_ _04665_ _04663_ _04664_ CPU.writeBack VGND VGND VPWR VPWR _05669_ sky130_fd_sc_hd__or4b_4
XFILLER_0_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10072_ _04666_ _05631_ VGND VGND VPWR VPWR _05632_ sky130_fd_sc_hd__nor2_2
XFILLER_0_100_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13900_ CPU.registerFile\[8\]\[30\] CPU.registerFile\[12\]\[30\] _07785_ VGND VGND
+ VPWR VPWR _08313_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_145_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783__231 clknet_1_1__leaf__07226_ VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__inv_2
X_13831_ _07370_ _08245_ VGND VGND VPWR VPWR _08246_ sky130_fd_sc_hd__or2_1
Xclkbuf_1_0__f__08433_ clknet_0__08433_ VGND VGND VPWR VPWR clknet_1_0__leaf__08433_
+ sky130_fd_sc_hd__clkbuf_16
X_13762_ CPU.registerFile\[3\]\[26\] _07373_ _07376_ VGND VGND VPWR VPWR _08179_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_39_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10974_ _06188_ VGND VGND VPWR VPWR _02021_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_48_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14425__556 clknet_1_0__leaf__02658_ VGND VGND VPWR VPWR net588 sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__08364_ clknet_0__08364_ VGND VGND VPWR VPWR clknet_1_0__leaf__08364_
+ sky130_fd_sc_hd__clkbuf_16
X_15501_ CPU.registerFile\[14\]\[4\] CPU.registerFile\[10\]\[4\] _02849_ VGND VGND
+ VPWR VPWR _02996_ sky130_fd_sc_hd__mux2_1
X_12713_ _07194_ VGND VGND VPWR VPWR _07195_ sky130_fd_sc_hd__buf_2
X_16481_ CPU.registerFile\[13\]\[31\] _02775_ VGND VGND VPWR VPWR _03949_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13693_ CPU.registerFile\[6\]\[24\] CPU.registerFile\[7\]\[24\] _07641_ VGND VGND
+ VPWR VPWR _08112_ sky130_fd_sc_hd__mux2_1
X_18220_ net61 _02500_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_15432_ CPU.registerFile\[25\]\[2\] _02928_ _02860_ VGND VGND VPWR VPWR _02929_ sky130_fd_sc_hd__o21a_1
X_12644_ net2313 _07146_ VGND VGND VPWR VPWR _00016_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_61_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18151_ clknet_leaf_28_clk _02431_ VGND VGND VPWR VPWR CPU.aluIn1\[17\] sky130_fd_sc_hd__dfxtp_4
X_12575_ CPU.registerFile\[4\]\[8\] _05252_ _07107_ VGND VGND VPWR VPWR _07111_ sky130_fd_sc_hd__mux2_1
X_15363_ _05405_ VGND VGND VPWR VPWR _02861_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17102_ _00012_ _00014_ VGND VGND VPWR VPWR CPU.mem_rstrb sky130_fd_sc_hd__dlxtn_2
XFILLER_0_81_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11526_ mapped_spi_ram.state\[2\] mapped_spi_ram.state\[1\] _06487_ VGND VGND VPWR
+ VPWR _06488_ sky130_fd_sc_hd__o21ai_1
X_18082_ net145 _02362_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15294_ CPU.registerFile\[24\]\[0\] _02789_ _02790_ _02792_ VGND VGND VPWR VPWR _02793_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_53_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17033_ net291 _01355_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_11457_ _06445_ VGND VGND VPWR VPWR _01795_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0__02722_ _02722_ VGND VGND VPWR VPWR clknet_0__02722_ sky130_fd_sc_hd__clkbuf_16
X_10408_ mapped_spi_flash.cmd_addr\[27\] _05825_ _05827_ mapped_spi_flash.cmd_addr\[28\]
+ VGND VGND VPWR VPWR _05835_ sky130_fd_sc_hd__a22o_1
X_14176_ _08425_ VGND VGND VPWR VPWR _01488_ sky130_fd_sc_hd__clkbuf_1
X_11388_ _05511_ net2009 _06408_ VGND VGND VPWR VPWR _06409_ sky130_fd_sc_hd__mux2_1
X_14471__598 clknet_1_1__leaf__02662_ VGND VGND VPWR VPWR net630 sky130_fd_sc_hd__inv_2
Xclkbuf_0__02653_ _02653_ VGND VGND VPWR VPWR clknet_0__02653_ sky130_fd_sc_hd__clkbuf_16
X_13127_ _07555_ _07560_ _07561_ _07563_ _07302_ VGND VGND VPWR VPWR _07564_ sky130_fd_sc_hd__a221o_1
X_10339_ _05516_ net2312 _05788_ VGND VGND VPWR VPWR _05791_ sky130_fd_sc_hd__mux2_1
X_13058_ _07397_ _07486_ _07496_ _07424_ VGND VGND VPWR VPWR _07497_ sky130_fd_sc_hd__a31o_1
X_17935_ net1124 _02219_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[15\] sky130_fd_sc_hd__dfxtp_1
X_12009_ _06773_ VGND VGND VPWR VPWR _01568_ sky130_fd_sc_hd__clkbuf_1
X_17866_ net1055 _02150_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_16817_ _07195_ _04117_ VGND VGND VPWR VPWR _04121_ sky130_fd_sc_hd__nor2_1
X_17797_ net986 _02081_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_14246__419 clknet_1_1__leaf__08434_ VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_37_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16748_ _04032_ CPU.PC\[15\] VGND VGND VPWR VPWR _04066_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16679_ _03995_ _05353_ _07123_ VGND VGND VPWR VPWR _04008_ sky130_fd_sc_hd__o21ai_1
X_09220_ _04811_ _04813_ _04815_ _04931_ VGND VGND VPWR VPWR _04932_ sky130_fd_sc_hd__or4b_4
XFILLER_0_72_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09151_ CPU.Bimm\[6\] _04819_ CPU.PC\[6\] VGND VGND VPWR VPWR _04863_ sky130_fd_sc_hd__a21oi_1
X_18349_ clknet_leaf_1_clk _02629_ VGND VGND VPWR VPWR per_uart.uart0.rx_count16\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09082_ _04350_ _04489_ _04792_ _04794_ VGND VGND VPWR VPWR _04795_ sky130_fd_sc_hd__a211o_1
XFILLER_0_32_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold800 CPU.registerFile\[18\]\[26\] VGND VGND VPWR VPWR net2041 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__03969_ _03969_ VGND VGND VPWR VPWR clknet_0__03969_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold811 CPU.registerFile\[26\]\[11\] VGND VGND VPWR VPWR net2052 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold822 CPU.registerFile\[18\]\[5\] VGND VGND VPWR VPWR net2063 sky130_fd_sc_hd__dlygate4sd3_1
Xhold833 CPU.registerFile\[17\]\[29\] VGND VGND VPWR VPWR net2074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 CPU.registerFile\[18\]\[1\] VGND VGND VPWR VPWR net2085 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold855 CPU.registerFile\[31\]\[28\] VGND VGND VPWR VPWR net2096 sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 CPU.registerFile\[1\]\[22\] VGND VGND VPWR VPWR net2107 sky130_fd_sc_hd__dlygate4sd3_1
X_14866__953 clknet_1_0__leaf__02702_ VGND VGND VPWR VPWR net985 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_92_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold877 CPU.registerFile\[20\]\[28\] VGND VGND VPWR VPWR net2118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 CPU.registerFile\[28\]\[15\] VGND VGND VPWR VPWR net2129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold899 CPU.registerFile\[7\]\[26\] VGND VGND VPWR VPWR net2140 sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ _05539_ net1903 _05581_ VGND VGND VPWR VPWR _05585_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__08358_ _08358_ VGND VGND VPWR VPWR clknet_0__08358_ sky130_fd_sc_hd__clkbuf_16
X_08935_ _04652_ _04216_ _04654_ VGND VGND VPWR VPWR _04655_ sky130_fd_sc_hd__a21o_1
X_08866_ CPU.state\[2\] CPU.state\[3\] net2 VGND VGND VPWR VPWR _04586_ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08797_ CPU.Iimm\[4\] CPU.Bimm\[4\] CPU.instr\[5\] VGND VGND VPWR VPWR _04517_ sky130_fd_sc_hd__mux2_4
Xclkbuf_1_0__f__02711_ clknet_0__02711_ VGND VGND VPWR VPWR clknet_1_0__leaf__02711_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_74_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_123_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09418_ _05118_ _05120_ _04373_ VGND VGND VPWR VPWR _05121_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10690_ _05497_ net2275 _06034_ VGND VGND VPWR VPWR _06038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09349_ net1242 _04442_ VGND VGND VPWR VPWR _05055_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_43_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12360_ _05150_ net1888 _06988_ VGND VGND VPWR VPWR _06997_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11311_ _06367_ VGND VGND VPWR VPWR _01863_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12291_ CPU.aluReg\[7\] _06953_ _06924_ VGND VGND VPWR VPWR _06954_ sky130_fd_sc_hd__mux2_1
X_11242_ net1606 _05683_ _06324_ VGND VGND VPWR VPWR _06331_ sky130_fd_sc_hd__mux2_1
X_11173_ _06294_ VGND VGND VPWR VPWR _01928_ sky130_fd_sc_hd__clkbuf_1
X_10124_ net2213 _05273_ _05655_ VGND VGND VPWR VPWR _05660_ sky130_fd_sc_hd__mux2_1
X_15981_ CPU.aluIn1\[16\] _03081_ _03463_ _03080_ VGND VGND VPWR VPWR _02430_ sky130_fd_sc_hd__o211a_1
X_17720_ net909 _02004_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_10055_ net1900 _05273_ _05618_ VGND VGND VPWR VPWR _05623_ sky130_fd_sc_hd__mux2_1
X_17651_ net840 _01939_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16602_ per_uart.uart0.rx_count16\[3\] per_uart.uart0.rx_count16\[2\] per_uart.uart0.rx_count16\[1\]
+ per_uart.uart0.rx_count16\[0\] VGND VGND VPWR VPWR _03973_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_3_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13814_ CPU.registerFile\[28\]\[27\] CPU.registerFile\[24\]\[27\] _07352_ VGND VGND
+ VPWR VPWR _08230_ sky130_fd_sc_hd__mux2_1
X_17582_ net771 _01870_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_34_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16533_ clknet_1_0__leaf__07219_ VGND VGND VPWR VPWR _03965_ sky130_fd_sc_hd__buf_1
X_13745_ CPU.registerFile\[31\]\[25\] _07482_ _07420_ CPU.registerFile\[27\]\[25\]
+ _07305_ VGND VGND VPWR VPWR _08163_ sky130_fd_sc_hd__o221a_1
X_10957_ net1577 _05668_ _06179_ VGND VGND VPWR VPWR _06180_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16464_ CPU.registerFile\[2\]\[31\] _03227_ _02873_ CPU.registerFile\[3\]\[31\] _03931_
+ VGND VGND VPWR VPWR _03932_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_158_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13676_ CPU.registerFile\[6\]\[23\] CPU.registerFile\[7\]\[23\] _07371_ VGND VGND
+ VPWR VPWR _08096_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_158_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10888_ _06142_ VGND VGND VPWR VPWR _06143_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_158_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18203_ net44 _02483_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15415_ CPU.registerFile\[15\]\[2\] _02826_ VGND VGND VPWR VPWR _02912_ sky130_fd_sc_hd__or2_1
XFILLER_0_26_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12627_ CPU.cycles\[3\] _07136_ VGND VGND VPWR VPWR _07138_ sky130_fd_sc_hd__and2_1
X_16395_ CPU.registerFile\[6\]\[29\] _02828_ VGND VGND VPWR VPWR _03865_ sky130_fd_sc_hd__or2_1
X_18134_ clknet_leaf_22_clk _02414_ VGND VGND VPWR VPWR CPU.aluIn1\[0\] sky130_fd_sc_hd__dfxtp_2
X_15346_ _02825_ _02842_ _02844_ VGND VGND VPWR VPWR _02845_ sky130_fd_sc_hd__o21a_1
XFILLER_0_26_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12558_ net2307 _05089_ _07096_ VGND VGND VPWR VPWR _07102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18065_ net1238 _02345_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_11509_ _06030_ _06475_ VGND VGND VPWR VPWR _01773_ sky130_fd_sc_hd__nor2_1
X_15277_ CPU.registerFile\[13\]\[0\] _02775_ VGND VGND VPWR VPWR _02776_ sky130_fd_sc_hd__or2_1
Xhold107 per_uart.uart0.enable16_counter\[9\] VGND VGND VPWR VPWR net1348 sky130_fd_sc_hd__dlygate4sd3_1
X_12489_ _07065_ VGND VGND VPWR VPWR _01345_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold118 mapped_spi_ram.cmd_addr\[9\] VGND VGND VPWR VPWR net1359 sky130_fd_sc_hd__dlygate4sd3_1
X_17016_ net274 _01338_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[10\] sky130_fd_sc_hd__dfxtp_1
Xhold129 mapped_spi_ram.cmd_addr\[18\] VGND VGND VPWR VPWR net1370 sky130_fd_sc_hd__dlygate4sd3_1
X_14588__703 clknet_1_0__leaf__02674_ VGND VGND VPWR VPWR net735 sky130_fd_sc_hd__inv_2
XFILLER_0_1_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__02705_ _02705_ VGND VGND VPWR VPWR clknet_0__02705_ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_74_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14159_ _08416_ VGND VGND VPWR VPWR _01480_ sky130_fd_sc_hd__clkbuf_1
X_14999__1073 clknet_1_1__leaf__02715_ VGND VGND VPWR VPWR net1105 sky130_fd_sc_hd__inv_2
XFILLER_0_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08720_ _04394_ _04438_ _04439_ VGND VGND VPWR VPWR _04440_ sky130_fd_sc_hd__o21a_1
X_17918_ net1107 _02202_ VGND VGND VPWR VPWR mapped_spi_flash.snd_bitcount\[4\] sky130_fd_sc_hd__dfxtp_1
X_08651_ _04222_ _04368_ _04370_ VGND VGND VPWR VPWR _04371_ sky130_fd_sc_hd__a21oi_1
X_17849_ net1038 _02133_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_14408__540 clknet_1_0__leaf__02657_ VGND VGND VPWR VPWR net572 sky130_fd_sc_hd__inv_2
X_08582_ CPU.mem_wdata\[0\] _04203_ _04301_ VGND VGND VPWR VPWR _04302_ sky130_fd_sc_hd__o21a_4
XFILLER_0_88_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_105_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_812 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09203_ _04499_ _04914_ VGND VGND VPWR VPWR _04915_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09134_ CPU.Jimm\[14\] _04829_ _04831_ VGND VGND VPWR VPWR _04846_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09065_ _04774_ _04775_ _04778_ VGND VGND VPWR VPWR _04779_ sky130_fd_sc_hd__or3_4
XFILLER_0_130_734 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold630 CPU.registerFile\[31\]\[8\] VGND VGND VPWR VPWR net1871 sky130_fd_sc_hd__dlygate4sd3_1
X_14454__582 clknet_1_0__leaf__02661_ VGND VGND VPWR VPWR net614 sky130_fd_sc_hd__inv_2
Xhold641 CPU.registerFile\[7\]\[24\] VGND VGND VPWR VPWR net1882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 CPU.registerFile\[29\]\[7\] VGND VGND VPWR VPWR net1893 sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 CPU.registerFile\[12\]\[2\] VGND VGND VPWR VPWR net1904 sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 CPU.registerFile\[13\]\[30\] VGND VGND VPWR VPWR net1915 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14192__370 clknet_1_1__leaf__08429_ VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__inv_2
Xhold685 CPU.registerFile\[26\]\[8\] VGND VGND VPWR VPWR net1926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 CPU.registerFile\[29\]\[2\] VGND VGND VPWR VPWR net1937 sky130_fd_sc_hd__dlygate4sd3_1
X_09967_ _05522_ net1714 _05570_ VGND VGND VPWR VPWR _05576_ sky130_fd_sc_hd__mux2_1
X_08918_ _04528_ net1280 _04506_ VGND VGND VPWR VPWR _04638_ sky130_fd_sc_hd__a21oi_1
X_09898_ _05532_ net1832 _05533_ VGND VGND VPWR VPWR _05534_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_125_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08849_ CPU.aluIn1\[17\] CPU.aluIn1\[16\] _04495_ VGND VGND VPWR VPWR _04569_ sky130_fd_sc_hd__o21ai_1
X_11860_ _06694_ VGND VGND VPWR VPWR _01638_ sky130_fd_sc_hd__clkbuf_1
X_10811_ _06101_ VGND VGND VPWR VPWR _02097_ sky130_fd_sc_hd__clkbuf_1
X_11791_ _05130_ net2243 _06650_ VGND VGND VPWR VPWR _06658_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_916 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13530_ CPU.registerFile\[18\]\[19\] CPU.registerFile\[22\]\[19\] _07457_ VGND VGND
+ VPWR VPWR _07954_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10742_ _05549_ CPU.registerFile\[28\]\[3\] _06056_ VGND VGND VPWR VPWR _06065_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13461_ CPU.registerFile\[9\]\[16\] _07619_ _07887_ VGND VGND VPWR VPWR _07888_ sky130_fd_sc_hd__o21a_1
X_10673_ net1357 _06018_ _06022_ _06027_ VGND VGND VPWR VPWR _02161_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_843 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12412_ _04982_ net2316 _07024_ VGND VGND VPWR VPWR _07025_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16180_ _03652_ _03653_ _03656_ _08401_ _02949_ VGND VGND VPWR VPWR _03657_ sky130_fd_sc_hd__a221o_1
X_13392_ CPU.registerFile\[15\]\[14\] _07276_ _07277_ CPU.registerFile\[11\]\[14\]
+ _07820_ VGND VGND VPWR VPWR _07821_ sky130_fd_sc_hd__o221a_1
XFILLER_0_63_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14537__657 clknet_1_0__leaf__02669_ VGND VGND VPWR VPWR net689 sky130_fd_sc_hd__inv_2
XFILLER_0_50_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_153_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12343_ _06976_ VGND VGND VPWR VPWR _06988_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_153_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12274_ CPU.aluIn1\[11\] _06940_ _06927_ VGND VGND VPWR VPWR _06941_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11225_ _06321_ VGND VGND VPWR VPWR _01903_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_56_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11156_ CPU.registerFile\[8\]\[1\] _05733_ _06251_ VGND VGND VPWR VPWR _06285_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10107_ net1898 _05109_ _05644_ VGND VGND VPWR VPWR _05651_ sky130_fd_sc_hd__mux2_1
X_11087_ net1858 _05733_ _06214_ VGND VGND VPWR VPWR _06248_ sky130_fd_sc_hd__mux2_1
X_15964_ _02885_ _03444_ _03445_ _03446_ _03054_ VGND VGND VPWR VPWR _03447_ sky130_fd_sc_hd__a221o_1
X_17703_ net892 _01991_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_10038_ net2278 _05109_ _05607_ VGND VGND VPWR VPWR _05614_ sky130_fd_sc_hd__mux2_1
X_15895_ CPU.registerFile\[29\]\[14\] _02800_ VGND VGND VPWR VPWR _03380_ sky130_fd_sc_hd__or2_1
X_14583__699 clknet_1_1__leaf__02673_ VGND VGND VPWR VPWR net731 sky130_fd_sc_hd__inv_2
X_17634_ net823 _01922_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17565_ net754 _01853_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_11989_ _05066_ net1884 _06758_ VGND VGND VPWR VPWR _06763_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13728_ CPU.registerFile\[21\]\[25\] _07265_ VGND VGND VPWR VPWR _08146_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17496_ net685 _01784_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16447_ CPU.registerFile\[31\]\[30\] _02887_ VGND VGND VPWR VPWR _03916_ sky130_fd_sc_hd__and2_1
X_13659_ net1530 _08018_ _08079_ _08017_ VGND VGND VPWR VPWR _01317_ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_140_Right_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16378_ CPU.registerFile\[1\]\[28\] _02814_ _03848_ _02816_ VGND VGND VPWR VPWR _03849_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18117_ net180 _02397_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15329_ _08394_ VGND VGND VPWR VPWR _02828_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18048_ net1221 _02328_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_09821_ net1927 _05359_ _05474_ VGND VGND VPWR VPWR _05482_ sky130_fd_sc_hd__mux2_1
X_09752_ _05440_ VGND VGND VPWR VPWR _05441_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_107_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08703_ _04406_ _04422_ _04277_ VGND VGND VPWR VPWR _04423_ sky130_fd_sc_hd__o21a_1
X_09683_ CPU.PC\[3\] CPU.PC\[2\] VGND VGND VPWR VPWR _05375_ sky130_fd_sc_hd__xnor2_1
X_08634_ _04351_ _04236_ _04353_ VGND VGND VPWR VPWR _04354_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_49_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ CPU.aluIn1\[4\] _04284_ VGND VGND VPWR VPWR _04285_ sky130_fd_sc_hd__or2_4
XFILLER_0_49_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08496_ _04215_ VGND VGND VPWR VPWR _04216_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_119_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_70_Left_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09117_ _04499_ _04292_ VGND VGND VPWR VPWR _04829_ sky130_fd_sc_hd__or2_2
XFILLER_0_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09048_ net1616 _04762_ _04668_ VGND VGND VPWR VPWR _04763_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold460 CPU.registerFile\[5\]\[19\] VGND VGND VPWR VPWR net1701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold471 CPU.registerFile\[7\]\[15\] VGND VGND VPWR VPWR net1712 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ _06207_ VGND VGND VPWR VPWR _02004_ sky130_fd_sc_hd__clkbuf_1
Xhold482 CPU.registerFile\[18\]\[22\] VGND VGND VPWR VPWR net1723 sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 CPU.registerFile\[29\]\[12\] VGND VGND VPWR VPWR net1734 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ _07234_ VGND VGND VPWR VPWR _07402_ sky130_fd_sc_hd__buf_4
Xhold1160 CPU.registerFile\[15\]\[8\] VGND VGND VPWR VPWR net2401 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1171 CPU.registerFile\[4\]\[12\] VGND VGND VPWR VPWR net2412 sky130_fd_sc_hd__dlygate4sd3_1
X_11912_ _06710_ VGND VGND VPWR VPWR _06722_ sky130_fd_sc_hd__clkbuf_4
Xhold1182 CPU.registerFile\[25\]\[12\] VGND VGND VPWR VPWR net2423 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15680_ _02786_ _03168_ _03170_ _02794_ VGND VGND VPWR VPWR _03171_ sky130_fd_sc_hd__a211o_1
X_12892_ _05232_ VGND VGND VPWR VPWR _07334_ sky130_fd_sc_hd__clkbuf_4
Xhold1193 CPU.registerFile\[29\]\[9\] VGND VGND VPWR VPWR net2434 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_300 _07320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_311 _07914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_322 _07914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_333 CPU.rs2\[25\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11843_ _06685_ VGND VGND VPWR VPWR _01646_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_344 _05338_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_355 _07268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_366 _02889_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17350_ net539 _01638_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[14\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_377 _07291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_388 _07271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14562_ clknet_1_0__leaf__02664_ VGND VGND VPWR VPWR _02672_ sky130_fd_sc_hd__buf_1
X_11774_ _04958_ net2204 _06639_ VGND VGND VPWR VPWR _06649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_399 _07250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16301_ CPU.registerFile\[6\]\[26\] CPU.registerFile\[7\]\[26\] _02870_ VGND VGND
+ VPWR VPWR _03774_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_155_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13513_ _07930_ _07937_ _07395_ VGND VGND VPWR VPWR _07938_ sky130_fd_sc_hd__o21a_1
X_14998__1072 clknet_1_1__leaf__02715_ VGND VGND VPWR VPWR net1104 sky130_fd_sc_hd__inv_2
X_17281_ net470 _01569_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10725_ _06033_ VGND VGND VPWR VPWR _06056_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_153_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_109_Left_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16232_ CPU.registerFile\[30\]\[24\] CPU.registerFile\[26\]\[24\] _03247_ VGND VGND
+ VPWR VPWR _03707_ sky130_fd_sc_hd__mux2_1
X_13444_ CPU.registerFile\[5\]\[16\] CPU.registerFile\[4\]\[16\] _07577_ VGND VGND
+ VPWR VPWR _07871_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10656_ _05817_ _05819_ VGND VGND VPWR VPWR _06014_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16163_ _08397_ _03635_ _03637_ _03639_ VGND VGND VPWR VPWR _03640_ sky130_fd_sc_hd__o22a_1
Xclkload16 clknet_leaf_20_clk VGND VGND VPWR VPWR clkload16/Y sky130_fd_sc_hd__clkinv_4
X_13375_ _04986_ VGND VGND VPWR VPWR _07804_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload27 clknet_leaf_11_clk VGND VGND VPWR VPWR clkload27/X sky130_fd_sc_hd__clkbuf_4
X_10587_ mapped_spi_flash.rcv_data\[27\] _05970_ VGND VGND VPWR VPWR _05975_ sky130_fd_sc_hd__or2_1
Xclkload38 clknet_1_0__leaf__02747_ VGND VGND VPWR VPWR clkload38/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_58_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload49 clknet_1_0__leaf__02715_ VGND VGND VPWR VPWR clkload49/Y sky130_fd_sc_hd__clkinvlp_4
X_12326_ _06979_ VGND VGND VPWR VPWR _01422_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16094_ CPU.registerFile\[20\]\[20\] _02855_ _03026_ VGND VGND VPWR VPWR _03573_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12257_ CPU.aluIn1\[15\] _06926_ _06927_ VGND VGND VPWR VPWR _06928_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11208_ _05537_ net2446 _06310_ VGND VGND VPWR VPWR _06313_ sky130_fd_sc_hd__mux2_1
X_12188_ CPU.aluIn1\[31\] _06874_ _06865_ VGND VGND VPWR VPWR _06875_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_118_Left_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11139_ _06276_ VGND VGND VPWR VPWR _01944_ sky130_fd_sc_hd__clkbuf_1
X_16996_ clknet_leaf_21_clk _01322_ VGND VGND VPWR VPWR CPU.rs2\[27\] sky130_fd_sc_hd__dfxtp_1
X_15947_ CPU.aluIn1\[15\] _02958_ _03413_ _03430_ _02995_ VGND VGND VPWR VPWR _02429_
+ sky130_fd_sc_hd__o221a_1
X_15878_ _02936_ _03356_ _03363_ _02934_ VGND VGND VPWR VPWR _03364_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_69_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17617_ net806 _01905_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_14829_ clknet_1_0__leaf__02697_ VGND VGND VPWR VPWR _02699_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_69_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17548_ net737 _01836_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_127_Left_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17479_ net668 net25 VGND VGND VPWR VPWR mapped_spi_flash.div_counter\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_82_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_136_Left_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09804_ net2105 _05170_ _05463_ VGND VGND VPWR VPWR _05473_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_89_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09735_ _05410_ _05414_ _05424_ VGND VGND VPWR VPWR _05425_ sky130_fd_sc_hd__or3_4
X_14566__683 clknet_1_1__leaf__02672_ VGND VGND VPWR VPWR net715 sky130_fd_sc_hd__inv_2
X_09666_ _05358_ VGND VGND VPWR VPWR _05359_ sky130_fd_sc_hd__buf_4
X_08617_ CPU.aluIn1\[18\] _04249_ VGND VGND VPWR VPWR _04337_ sky130_fd_sc_hd__nand2_1
X_09597_ _05291_ _04918_ VGND VGND VPWR VPWR _05292_ sky130_fd_sc_hd__xnor2_1
X_08548_ CPU.rs2\[9\] CPU.Bimm\[9\] net1296 VGND VGND VPWR VPWR _04268_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_137_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08479_ _04196_ _04197_ _04198_ VGND VGND VPWR VPWR _04199_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_64_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10510_ _04539_ _05915_ VGND VGND VPWR VPWR _05916_ sky130_fd_sc_hd__or2_1
X_11490_ _06462_ VGND VGND VPWR VPWR _01779_ sky130_fd_sc_hd__clkbuf_1
X_18372__31 VGND VGND VPWR VPWR _18372__31/HI net31 sky130_fd_sc_hd__conb_1
XFILLER_0_134_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10441_ _05852_ _04608_ VGND VGND VPWR VPWR _05859_ sky130_fd_sc_hd__nor2_1
X_14731__831 clknet_1_1__leaf__02689_ VGND VGND VPWR VPWR net863 sky130_fd_sc_hd__inv_2
XFILLER_0_150_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_150_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_150_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13160_ _07412_ _07594_ _07595_ VGND VGND VPWR VPWR _07596_ sky130_fd_sc_hd__o21a_1
X_10372_ _05549_ net2287 _05799_ VGND VGND VPWR VPWR _05808_ sky130_fd_sc_hd__mux2_1
X_12111_ _06827_ VGND VGND VPWR VPWR _01519_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13091_ _07351_ _07528_ VGND VGND VPWR VPWR _07529_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_53_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12042_ _04798_ net1866 _06783_ VGND VGND VPWR VPWR _06791_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_53_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14649__758 clknet_1_0__leaf__02680_ VGND VGND VPWR VPWR net790 sky130_fd_sc_hd__inv_2
Xhold290 CPU.rs2\[27\] VGND VGND VPWR VPWR net1531 sky130_fd_sc_hd__dlygate4sd3_1
X_16850_ net1553 VGND VGND VPWR VPWR _02619_ sky130_fd_sc_hd__clkbuf_1
X_15801_ _03285_ _03286_ _03288_ _02945_ VGND VGND VPWR VPWR _03289_ sky130_fd_sc_hd__o22a_2
XTAP_TAPCELL_ROW_148_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16781_ _05289_ _04995_ _07132_ VGND VGND VPWR VPWR _04094_ sky130_fd_sc_hd__o21ai_1
X_15732_ _03030_ _03220_ _03221_ _02901_ VGND VGND VPWR VPWR _03222_ sky130_fd_sc_hd__a22o_1
X_12944_ _07364_ _07384_ VGND VGND VPWR VPWR _07385_ sky130_fd_sc_hd__or2_1
X_15663_ _03072_ _03153_ _03154_ VGND VGND VPWR VPWR _03155_ sky130_fd_sc_hd__o21a_1
XANTENNA_130 _05545_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12875_ CPU.registerFile\[5\]\[1\] CPU.registerFile\[4\]\[1\] net14 VGND VGND VPWR
+ VPWR _07317_ sky130_fd_sc_hd__mux2_1
XANTENNA_141 _05710_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_152 _07271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17402_ net591 _01690_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_bitcount\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11826_ net1627 _05673_ _06675_ VGND VGND VPWR VPWR _06677_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_163 _07322_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15594_ CPU.registerFile\[15\]\[6\] CPU.registerFile\[11\]\[6\] _02773_ VGND VGND
+ VPWR VPWR _03087_ sky130_fd_sc_hd__mux2_1
XANTENNA_174 _07476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_185 _07744_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_196 _07841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17333_ net522 _01621_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11757_ _06640_ VGND VGND VPWR VPWR _01687_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__03971_ clknet_0__03971_ VGND VGND VPWR VPWR clknet_1_1__leaf__03971_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_64_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14023__302 clknet_1_0__leaf__08362_ VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__inv_2
XFILLER_0_138_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10708_ _06047_ VGND VGND VPWR VPWR _02146_ sky130_fd_sc_hd__clkbuf_1
X_17264_ net454 _01552_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_14394__528 clknet_1_0__leaf__02655_ VGND VGND VPWR VPWR net560 sky130_fd_sc_hd__inv_2
XFILLER_0_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11688_ net1424 _06588_ VGND VGND VPWR VPWR _06597_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16215_ _03689_ _03690_ _08400_ VGND VGND VPWR VPWR _03691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload105 clknet_1_1__leaf__08360_ VGND VGND VPWR VPWR clkload105/Y sky130_fd_sc_hd__clkinvlp_4
X_13427_ CPU.registerFile\[28\]\[15\] CPU.registerFile\[24\]\[15\] _07292_ VGND VGND
+ VPWR VPWR _07855_ sky130_fd_sc_hd__mux2_1
Xclkload116 clknet_1_0__leaf__03966_ VGND VGND VPWR VPWR clkload116/Y sky130_fd_sc_hd__clkinvlp_4
X_17195_ clknet_leaf_11_clk _01483_ VGND VGND VPWR VPWR CPU.Bimm\[5\] sky130_fd_sc_hd__dfxtp_2
X_10639_ net1486 _05994_ VGND VGND VPWR VPWR _06004_ sky130_fd_sc_hd__or2_1
XFILLER_0_141_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16146_ CPU.registerFile\[16\]\[21\] _02831_ _02834_ CPU.registerFile\[17\]\[21\]
+ _02854_ VGND VGND VPWR VPWR _03624_ sky130_fd_sc_hd__o221a_1
XFILLER_0_11_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__08360_ clknet_0__08360_ VGND VGND VPWR VPWR clknet_1_1__leaf__08360_
+ sky130_fd_sc_hd__clkbuf_16
X_13358_ _07273_ _07786_ _07787_ VGND VGND VPWR VPWR _07788_ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12309_ CPU.aluReg\[3\] CPU.aluReg\[1\] _06939_ VGND VGND VPWR VPWR _06967_ sky130_fd_sc_hd__mux2_1
X_16077_ CPU.registerFile\[27\]\[19\] _02928_ _02923_ VGND VGND VPWR VPWR _03557_
+ sky130_fd_sc_hd__o21a_1
X_13289_ _07713_ _07720_ _07395_ VGND VGND VPWR VPWR _07721_ sky130_fd_sc_hd__o21a_1
XFILLER_0_122_895 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15028_ clknet_1_1__leaf__02708_ VGND VGND VPWR VPWR _02718_ sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14860__948 clknet_1_1__leaf__02701_ VGND VGND VPWR VPWR net980 sky130_fd_sc_hd__inv_2
XFILLER_0_127_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput3 spi_miso VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_1
X_16979_ clknet_leaf_26_clk _01305_ VGND VGND VPWR VPWR CPU.rs2\[10\] sky130_fd_sc_hd__dfxtp_1
X_09520_ _05217_ _04428_ VGND VGND VPWR VPWR _05218_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_84_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09451_ mapped_spi_ram.rcv_data\[20\] _04689_ _04691_ mapped_spi_flash.rcv_data\[20\]
+ VGND VGND VPWR VPWR _05152_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09382_ _04925_ _05086_ VGND VGND VPWR VPWR _05087_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_144_Left_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14997__1071 clknet_1_1__leaf__02715_ VGND VGND VPWR VPWR net1103 sky130_fd_sc_hd__inv_2
X_09718_ mapped_spi_flash.rcv_data\[25\] _04784_ _05407_ VGND VGND VPWR VPWR _05408_
+ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_153_Left_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10990_ net1725 _05704_ _06190_ VGND VGND VPWR VPWR _06197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09649_ _05275_ _05335_ _05341_ _05286_ VGND VGND VPWR VPWR _05342_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_679 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16589__60 clknet_1_1__leaf__03970_ VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__inv_2
X_12660_ CPU.cycles\[16\] _07154_ net1416 VGND VGND VPWR VPWR _07157_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11611_ net1362 _06494_ _06544_ _06539_ VGND VGND VPWR VPWR _01736_ sky130_fd_sc_hd__o211a_1
X_12591_ net1641 _05447_ _07084_ VGND VGND VPWR VPWR _07119_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_705 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11542_ mapped_spi_ram.cmd_addr\[23\] _06493_ VGND VGND VPWR VPWR _06497_ sky130_fd_sc_hd__and2b_1
X_14261_ _05183_ _05201_ _05216_ _08439_ VGND VGND VPWR VPWR _08440_ sky130_fd_sc_hd__or4_1
XFILLER_0_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11473_ _06453_ VGND VGND VPWR VPWR _01787_ sky130_fd_sc_hd__clkbuf_1
X_16000_ _03195_ _03479_ _03480_ _03481_ _03245_ VGND VGND VPWR VPWR _03482_ sky130_fd_sc_hd__a221o_1
X_13212_ _07302_ VGND VGND VPWR VPWR _07646_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_122_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10424_ _05830_ _05845_ VGND VGND VPWR VPWR _05846_ sky130_fd_sc_hd__and2_1
XFILLER_0_61_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13143_ CPU.registerFile\[1\]\[7\] _07576_ _07578_ _07369_ VGND VGND VPWR VPWR _07579_
+ sky130_fd_sc_hd__a22o_1
X_10355_ _05776_ VGND VGND VPWR VPWR _05799_ sky130_fd_sc_hd__buf_4
X_13074_ CPU.registerFile\[1\]\[5\] _07255_ _07511_ _07318_ VGND VGND VPWR VPWR _07512_
+ sky130_fd_sc_hd__a22o_1
X_10286_ _05739_ VGND VGND VPWR VPWR _05762_ sky130_fd_sc_hd__buf_4
X_17951_ net1140 _02235_ VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dfxtp_1
X_12025_ _06781_ VGND VGND VPWR VPWR _01560_ sky130_fd_sc_hd__clkbuf_1
X_16902_ CPU.mem_wdata\[2\] _04174_ _04178_ _04176_ VGND VGND VPWR VPWR _02636_ sky130_fd_sc_hd__o211a_1
X_17882_ net1071 _02166_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[0\] sky130_fd_sc_hd__dfxtp_1
X_16833_ _04131_ _04132_ VGND VGND VPWR VPWR _04133_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16764_ _08457_ _04077_ _04078_ _04079_ VGND VGND VPWR VPWR _04080_ sky130_fd_sc_hd__a31oi_1
X_13976_ clknet_1_1__leaf__07223_ VGND VGND VPWR VPWR _08358_ sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15715_ _08405_ _03203_ _03204_ VGND VGND VPWR VPWR _03205_ sky130_fd_sc_hd__a21o_1
XFILLER_0_158_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12927_ _05284_ VGND VGND VPWR VPWR _07368_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_66_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16695_ _03991_ net1590 VGND VGND VPWR VPWR _04021_ sky130_fd_sc_hd__nand2_1
X_12760__210 clknet_1_1__leaf__07224_ VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15646_ _02809_ VGND VGND VPWR VPWR _03138_ sky130_fd_sc_hd__buf_4
X_12858_ CPU.registerFile\[29\]\[0\] _07289_ _07290_ CPU.registerFile\[25\]\[0\] _07300_
+ VGND VGND VPWR VPWR _07301_ sky130_fd_sc_hd__o221a_1
XFILLER_0_158_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14402__535 clknet_1_0__leaf__02656_ VGND VGND VPWR VPWR net567 sky130_fd_sc_hd__inv_2
X_11809_ _06667_ VGND VGND VPWR VPWR _01662_ sky130_fd_sc_hd__clkbuf_1
X_18365_ clknet_leaf_9_clk _02643_ VGND VGND VPWR VPWR per_uart.d_in_uart\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15577_ _03065_ _03067_ _03070_ VGND VGND VPWR VPWR _03071_ sky130_fd_sc_hd__o21a_1
X_12789_ _07231_ VGND VGND VPWR VPWR _07232_ sky130_fd_sc_hd__buf_4
X_17316_ net505 _01604_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18296_ net129 _02576_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17247_ net437 _01535_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17178_ clknet_leaf_25_clk _01466_ VGND VGND VPWR VPWR CPU.Bimm\[1\] sky130_fd_sc_hd__dfxtp_1
X_16129_ _03602_ _03606_ _08410_ VGND VGND VPWR VPWR _03607_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15184__1209 clknet_1_1__leaf__02748_ VGND VGND VPWR VPWR net1241 sky130_fd_sc_hd__inv_2
X_08951_ CPU.Bimm\[10\] _04372_ VGND VGND VPWR VPWR _04670_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_94_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__02698_ clknet_0__02698_ VGND VGND VPWR VPWR clknet_1_1__leaf__02698_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_138_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__07225_ clknet_0__07225_ VGND VGND VPWR VPWR clknet_1_1__leaf__07225_
+ sky130_fd_sc_hd__clkbuf_16
X_08882_ _04559_ _04562_ _04563_ VGND VGND VPWR VPWR _04602_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09503_ _04269_ _04318_ VGND VGND VPWR VPWR _05202_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_616 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09434_ _04850_ _04894_ VGND VGND VPWR VPWR _05136_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14678__784 clknet_1_0__leaf__02683_ VGND VGND VPWR VPWR net816 sky130_fd_sc_hd__inv_2
XFILLER_0_136_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09365_ _05069_ VGND VGND VPWR VPWR _05070_ sky130_fd_sc_hd__buf_4
X_14377__512 clknet_1_0__leaf__02654_ VGND VGND VPWR VPWR net544 sky130_fd_sc_hd__inv_2
XFILLER_0_90_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_30 _03064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09296_ _04928_ _05004_ VGND VGND VPWR VPWR _05005_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_10_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_41 _03728_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_52 _04957_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_63 _05046_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_74 _05149_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_85 _05253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_96 _05333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10140_ _04658_ VGND VGND VPWR VPWR _05668_ sky130_fd_sc_hd__clkbuf_4
X_10071_ _04661_ _04660_ VGND VGND VPWR VPWR _05631_ sky130_fd_sc_hd__nand2b_4
X_14843__932 clknet_1_1__leaf__02700_ VGND VGND VPWR VPWR net964 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_145_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13830_ CPU.registerFile\[30\]\[28\] CPU.registerFile\[26\]\[28\] _04936_ VGND VGND
+ VPWR VPWR _08245_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__08432_ clknet_0__08432_ VGND VGND VPWR VPWR clknet_1_0__leaf__08432_
+ sky130_fd_sc_hd__clkbuf_16
Xmax_cap21 _06485_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_1
X_13761_ CPU.registerFile\[2\]\[26\] _07322_ VGND VGND VPWR VPWR _08178_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_39_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10973_ net1680 _05687_ _06179_ VGND VGND VPWR VPWR _06188_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__08363_ clknet_0__08363_ VGND VGND VPWR VPWR clknet_1_0__leaf__08363_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15500_ CPU.aluIn1\[3\] _02958_ _02977_ _02994_ _02995_ VGND VGND VPWR VPWR _02417_
+ sky130_fd_sc_hd__o221a_1
X_12712_ per_uart.uart0.enable16_counter\[15\] _07193_ VGND VGND VPWR VPWR _07194_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_57_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16480_ CPU.registerFile\[9\]\[31\] _08404_ _02860_ VGND VGND VPWR VPWR _03948_ sky130_fd_sc_hd__o21a_1
X_13692_ CPU.rs2\[23\] _07705_ _08095_ _08111_ _07737_ VGND VGND VPWR VPWR _01318_
+ sky130_fd_sc_hd__o221a_1
X_15431_ _05406_ VGND VGND VPWR VPWR _02928_ sky130_fd_sc_hd__buf_4
X_12643_ _07146_ _07147_ VGND VGND VPWR VPWR _00046_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18150_ clknet_leaf_19_clk _02430_ VGND VGND VPWR VPWR CPU.aluIn1\[16\] sky130_fd_sc_hd__dfxtp_4
X_15362_ _05070_ VGND VGND VPWR VPWR _02860_ sky130_fd_sc_hd__clkbuf_4
X_12574_ _07110_ VGND VGND VPWR VPWR _01272_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_61_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_902 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17101_ net359 _01423_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11525_ _06471_ _06486_ VGND VGND VPWR VPWR _06487_ sky130_fd_sc_hd__nor2_1
X_18081_ net144 _02361_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_15293_ CPU.registerFile\[28\]\[0\] _02791_ VGND VGND VPWR VPWR _02792_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17032_ net290 _01354_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_11456_ _05511_ net2475 _06444_ VGND VGND VPWR VPWR _06445_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__02721_ _02721_ VGND VGND VPWR VPWR clknet_0__02721_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10407_ _05834_ VGND VGND VPWR VPWR _02233_ sky130_fd_sc_hd__clkbuf_1
X_14175_ CPU.Bimm\[10\] _04692_ _07127_ VGND VGND VPWR VPWR _08425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11387_ _06396_ VGND VGND VPWR VPWR _06408_ sky130_fd_sc_hd__buf_4
XFILLER_0_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__02652_ _02652_ VGND VGND VPWR VPWR clknet_0__02652_ sky130_fd_sc_hd__clkbuf_16
X_13126_ _07351_ _07562_ VGND VGND VPWR VPWR _07563_ sky130_fd_sc_hd__or2_1
X_10338_ _05790_ VGND VGND VPWR VPWR _02259_ sky130_fd_sc_hd__clkbuf_1
X_13057_ _07411_ _07491_ _07495_ VGND VGND VPWR VPWR _07496_ sky130_fd_sc_hd__or3_1
X_17934_ net1123 _02218_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[14\] sky130_fd_sc_hd__dfxtp_1
X_10269_ _05753_ VGND VGND VPWR VPWR _02306_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12008_ _05253_ net2108 _06769_ VGND VGND VPWR VPWR _06773_ sky130_fd_sc_hd__mux2_1
X_17865_ net1054 _02149_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_16816_ _04120_ VGND VGND VPWR VPWR _02608_ sky130_fd_sc_hd__clkbuf_1
X_17796_ net985 _02080_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_16747_ _04061_ _04065_ _04015_ VGND VGND VPWR VPWR _02594_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_17_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16678_ _08379_ _05347_ _04006_ VGND VGND VPWR VPWR _04007_ sky130_fd_sc_hd__or3b_1
XFILLER_0_119_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16568__41 clknet_1_1__leaf__03968_ VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__inv_2
X_15629_ _02759_ _03116_ _03120_ _02767_ VGND VGND VPWR VPWR _03121_ sky130_fd_sc_hd__a211o_1
XFILLER_0_57_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09150_ CPU.PC\[6\] CPU.Bimm\[6\] _04819_ VGND VGND VPWR VPWR _04862_ sky130_fd_sc_hd__and3_1
X_18348_ clknet_leaf_1_clk _02628_ VGND VGND VPWR VPWR per_uart.uart0.rx_count16\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14996__1070 clknet_1_0__leaf__02715_ VGND VGND VPWR VPWR net1102 sky130_fd_sc_hd__inv_2
XFILLER_0_71_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16583__55 clknet_1_0__leaf__03969_ VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__inv_2
X_09081_ _04236_ _04698_ _04218_ CPU.aluReg\[24\] _04793_ VGND VGND VPWR VPWR _04794_
+ sky130_fd_sc_hd__a221o_1
X_18279_ net112 _02559_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15227__137 clknet_1_0__leaf__02753_ VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__inv_2
XFILLER_0_141_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__03968_ _03968_ VGND VGND VPWR VPWR clknet_0__03968_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_140_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold801 CPU.registerFile\[15\]\[12\] VGND VGND VPWR VPWR net2042 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_730 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold812 CPU.registerFile\[24\]\[14\] VGND VGND VPWR VPWR net2053 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold823 mapped_spi_flash.rcv_data\[10\] VGND VGND VPWR VPWR net2064 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold834 CPU.registerFile\[3\]\[29\] VGND VGND VPWR VPWR net2075 sky130_fd_sc_hd__dlygate4sd3_1
Xhold845 CPU.registerFile\[29\]\[20\] VGND VGND VPWR VPWR net2086 sky130_fd_sc_hd__dlygate4sd3_1
X_14001__282 clknet_1_0__leaf__08360_ VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__inv_2
Xhold856 CPU.registerFile\[31\]\[25\] VGND VGND VPWR VPWR net2097 sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 CPU.registerFile\[12\]\[8\] VGND VGND VPWR VPWR net2108 sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 CPU.registerFile\[29\]\[30\] VGND VGND VPWR VPWR net2119 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09983_ _05584_ VGND VGND VPWR VPWR _02455_ sky130_fd_sc_hd__clkbuf_1
Xhold889 CPU.registerFile\[28\]\[5\] VGND VGND VPWR VPWR net2130 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__08357_ _08357_ VGND VGND VPWR VPWR clknet_0__08357_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08934_ _04372_ _04292_ _04653_ VGND VGND VPWR VPWR _04654_ sky130_fd_sc_hd__or3_4
X_08865_ _04577_ _04583_ _04579_ VGND VGND VPWR VPWR _04585_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_127_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__02710_ clknet_0__02710_ VGND VGND VPWR VPWR clknet_1_0__leaf__02710_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_98_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08796_ CPU.aluIn1\[7\] CPU.Bimm\[7\] VGND VGND VPWR VPWR _04516_ sky130_fd_sc_hd__or2_2
XPHY_EDGE_ROW_154_Right_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_140_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09417_ _04438_ _05119_ VGND VGND VPWR VPWR _05120_ sky130_fd_sc_hd__and2b_1
XFILLER_0_109_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09348_ _04443_ _05053_ VGND VGND VPWR VPWR _05054_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_43_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09279_ _04782_ _04987_ _04777_ VGND VGND VPWR VPWR _04988_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11310_ _05503_ net2345 _06360_ VGND VGND VPWR VPWR _06367_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12290_ CPU.aluIn1\[7\] _06952_ _06927_ VGND VGND VPWR VPWR _06953_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11241_ _06330_ VGND VGND VPWR VPWR _01896_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11172_ _05501_ net1645 _06288_ VGND VGND VPWR VPWR _06294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14431__561 clknet_1_1__leaf__02659_ VGND VGND VPWR VPWR net593 sky130_fd_sc_hd__inv_2
X_10123_ _05659_ VGND VGND VPWR VPWR _02358_ sky130_fd_sc_hd__clkbuf_1
X_15980_ _08407_ _03439_ _03448_ _03462_ _07424_ VGND VGND VPWR VPWR _03463_ sky130_fd_sc_hd__a311o_2
X_10054_ _05622_ VGND VGND VPWR VPWR _02390_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17650_ net839 _01938_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_14862_ clknet_1_0__leaf__02697_ VGND VGND VPWR VPWR _02702_ sky130_fd_sc_hd__buf_1
XFILLER_0_54_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14349__488 clknet_1_1__leaf__08467_ VGND VGND VPWR VPWR net520 sky130_fd_sc_hd__inv_2
X_16601_ per_uart.uart0.rx_busy VGND VGND VPWR VPWR _03972_ sky130_fd_sc_hd__inv_2
X_13813_ CPU.registerFile\[29\]\[27\] _07502_ _07348_ CPU.registerFile\[25\]\[27\]
+ _07300_ VGND VGND VPWR VPWR _08229_ sky130_fd_sc_hd__o221a_1
X_17581_ net770 _01869_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_3_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_121_Right_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13744_ CPU.registerFile\[30\]\[25\] CPU.registerFile\[26\]\[25\] _07492_ VGND VGND
+ VPWR VPWR _08162_ sky130_fd_sc_hd__mux2_1
X_10956_ _06178_ VGND VGND VPWR VPWR _06179_ sky130_fd_sc_hd__buf_4
X_14961__1039 clknet_1_1__leaf__02711_ VGND VGND VPWR VPWR net1071 sky130_fd_sc_hd__inv_2
XFILLER_0_85_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15183__1208 clknet_1_1__leaf__02748_ VGND VGND VPWR VPWR net1240 sky130_fd_sc_hd__inv_2
X_16463_ CPU.registerFile\[7\]\[31\] _02898_ _02999_ _03930_ VGND VGND VPWR VPWR _03931_
+ sky130_fd_sc_hd__o211a_1
X_13675_ _07394_ _08087_ _08091_ _08094_ _07232_ VGND VGND VPWR VPWR _08095_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_158_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10887_ _05594_ _06141_ VGND VGND VPWR VPWR _06142_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_158_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18202_ net43 _02482_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_15414_ _02910_ VGND VGND VPWR VPWR _02911_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_158_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12626_ _07136_ net1420 VGND VGND VPWR VPWR _00037_ sky130_fd_sc_hd__nor2_1
X_16394_ CPU.registerFile\[1\]\[29\] _03228_ _03863_ _02818_ VGND VGND VPWR VPWR _03864_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18133_ net196 _02413_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_15345_ _02843_ VGND VGND VPWR VPWR _02844_ sky130_fd_sc_hd__buf_4
X_12557_ _07101_ VGND VGND VPWR VPWR _01280_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18064_ net1237 _02344_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_11508_ net1516 _06473_ _06474_ VGND VGND VPWR VPWR _06475_ sky130_fd_sc_hd__a21oi_1
X_15276_ _02760_ VGND VGND VPWR VPWR _02775_ sky130_fd_sc_hd__clkbuf_4
X_12488_ net2054 _05700_ _07060_ VGND VGND VPWR VPWR _07065_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold108 mapped_spi_ram.rcv_bitcount\[2\] VGND VGND VPWR VPWR net1349 sky130_fd_sc_hd__dlygate4sd3_1
X_17015_ net273 _01337_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_14059__334 clknet_1_0__leaf__08366_ VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__inv_2
X_14514__636 clknet_1_0__leaf__02667_ VGND VGND VPWR VPWR net668 sky130_fd_sc_hd__inv_2
Xhold119 mapped_spi_flash.cmd_addr\[17\] VGND VGND VPWR VPWR net1360 sky130_fd_sc_hd__dlygate4sd3_1
X_11439_ _05495_ net2432 _06433_ VGND VGND VPWR VPWR _06436_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__02704_ _02704_ VGND VGND VPWR VPWR clknet_0__02704_ sky130_fd_sc_hd__clkbuf_16
X_14252__424 clknet_1_1__leaf__08435_ VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__inv_2
X_14158_ CPU.Iimm\[2\] _07369_ _08413_ VGND VGND VPWR VPWR _08416_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_74_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ _07254_ _07541_ _07545_ _07268_ VGND VGND VPWR VPWR _07546_ sky130_fd_sc_hd__o211a_1
X_14089_ _08370_ VGND VGND VPWR VPWR _01456_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17917_ net1106 _02201_ VGND VGND VPWR VPWR mapped_spi_flash.snd_bitcount\[3\] sky130_fd_sc_hd__dfxtp_1
X_08650_ _04369_ _04207_ VGND VGND VPWR VPWR _04370_ sky130_fd_sc_hd__xnor2_2
X_17848_ net1037 _02132_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_08581_ _04293_ _04294_ _04295_ _04291_ CPU.Iimm\[0\] VGND VGND VPWR VPWR _04301_
+ sky130_fd_sc_hd__a221o_1
X_17779_ net968 _02063_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_105_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14560__678 clknet_1_0__leaf__02671_ VGND VGND VPWR VPWR net710 sky130_fd_sc_hd__inv_2
XFILLER_0_49_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_105_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09202_ net1274 CPU.instr\[2\] _04291_ _04830_ VGND VGND VPWR VPWR _04914_ sky130_fd_sc_hd__and4_1
XFILLER_0_56_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09133_ CPU.PC\[15\] _04844_ VGND VGND VPWR VPWR _04845_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09064_ _04216_ _04776_ net1277 VGND VGND VPWR VPWR _04778_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_115_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold620 CPU.registerFile\[31\]\[18\] VGND VGND VPWR VPWR net1861 sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 CPU.registerFile\[7\]\[25\] VGND VGND VPWR VPWR net1872 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold642 CPU.registerFile\[23\]\[13\] VGND VGND VPWR VPWR net1883 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14489__613 clknet_1_0__leaf__02665_ VGND VGND VPWR VPWR net645 sky130_fd_sc_hd__inv_2
Xhold653 CPU.registerFile\[16\]\[7\] VGND VGND VPWR VPWR net1894 sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 CPU.registerFile\[3\]\[8\] VGND VGND VPWR VPWR net1905 sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 CPU.registerFile\[21\]\[2\] VGND VGND VPWR VPWR net1916 sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 CPU.registerFile\[19\]\[4\] VGND VGND VPWR VPWR net1927 sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 CPU.registerFile\[27\]\[6\] VGND VGND VPWR VPWR net1938 sky130_fd_sc_hd__dlygate4sd3_1
X_09966_ _05575_ VGND VGND VPWR VPWR _02463_ sky130_fd_sc_hd__clkbuf_1
X_08917_ _04624_ _04636_ VGND VGND VPWR VPWR _04637_ sky130_fd_sc_hd__nand2_1
X_09897_ _05490_ VGND VGND VPWR VPWR _05533_ sky130_fd_sc_hd__clkbuf_4
X_08848_ _04566_ _04567_ VGND VGND VPWR VPWR _04568_ sky130_fd_sc_hd__nand2_1
X_14229__404 clknet_1_0__leaf__08432_ VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__inv_2
X_08779_ CPU.instr\[3\] VGND VGND VPWR VPWR _04499_ sky130_fd_sc_hd__buf_2
XFILLER_0_68_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ _05549_ net1683 _06092_ VGND VGND VPWR VPWR _06101_ sky130_fd_sc_hd__mux2_1
X_11790_ _06657_ VGND VGND VPWR VPWR _01671_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10741_ _06064_ VGND VGND VPWR VPWR _02130_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13460_ CPU.registerFile\[13\]\[16\] _07629_ _07886_ _07371_ _04971_ VGND VGND VPWR
+ VPWR _07887_ sky130_fd_sc_hd__o221a_1
X_16547__22 clknet_1_1__leaf__03966_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__inv_2
XFILLER_0_48_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10672_ _05963_ _06026_ VGND VGND VPWR VPWR _06027_ sky130_fd_sc_hd__nand2_1
XFILLER_0_75_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12411_ _07012_ VGND VGND VPWR VPWR _07024_ sky130_fd_sc_hd__buf_4
XFILLER_0_152_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13391_ _07252_ VGND VGND VPWR VPWR _07820_ sky130_fd_sc_hd__buf_4
XFILLER_0_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_20_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_8
X_15130_ clknet_1_1__leaf__02720_ VGND VGND VPWR VPWR _02744_ sky130_fd_sc_hd__buf_1
X_16562__36 clknet_1_1__leaf__03967_ VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__inv_2
X_12342_ _06987_ VGND VGND VPWR VPWR _01414_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12273_ CPU.aluReg\[12\] CPU.aluReg\[10\] _06939_ VGND VGND VPWR VPWR _06940_ sky130_fd_sc_hd__mux2_1
X_11224_ _05553_ net2126 _06287_ VGND VGND VPWR VPWR _06321_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11155_ _06284_ VGND VGND VPWR VPWR _01936_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_8_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10106_ _05650_ VGND VGND VPWR VPWR _02366_ sky130_fd_sc_hd__clkbuf_1
X_11086_ _06247_ VGND VGND VPWR VPWR _01968_ sky130_fd_sc_hd__clkbuf_1
X_15963_ CPU.registerFile\[25\]\[16\] _03280_ _02940_ VGND VGND VPWR VPWR _03446_
+ sky130_fd_sc_hd__o21a_1
X_17702_ net891 _01990_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_10037_ _05613_ VGND VGND VPWR VPWR _02398_ sky130_fd_sc_hd__clkbuf_1
X_15894_ CPU.registerFile\[27\]\[14\] CPU.registerFile\[31\]\[14\] _03050_ VGND VGND
+ VPWR VPWR _03379_ sky130_fd_sc_hd__mux2_1
X_14702__806 clknet_1_0__leaf__02685_ VGND VGND VPWR VPWR net838 sky130_fd_sc_hd__inv_2
X_15256__163 clknet_1_1__leaf__02756_ VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__inv_2
X_17633_ net822 _01921_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_17564_ net753 _01852_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_11988_ _06762_ VGND VGND VPWR VPWR _01578_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13727_ _04814_ _08142_ _08144_ _04987_ VGND VGND VPWR VPWR _08145_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_27_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10939_ net1558 _05721_ _06165_ VGND VGND VPWR VPWR _06170_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_27_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17495_ net684 _01783_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13658_ _07394_ _08064_ _08078_ _08015_ VGND VGND VPWR VPWR _08079_ sky130_fd_sc_hd__a211o_1
X_16446_ CPU.registerFile\[25\]\[30\] CPU.registerFile\[29\]\[30\] _02798_ VGND VGND
+ VPWR VPWR _03915_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12609_ _07127_ VGND VGND VPWR VPWR _00000_ sky130_fd_sc_hd__clkbuf_4
X_16377_ CPU.registerFile\[5\]\[28\] CPU.registerFile\[4\]\[28\] _02805_ VGND VGND
+ VPWR VPWR _03848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13589_ _07330_ _08011_ VGND VGND VPWR VPWR _08012_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_11_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_30_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15328_ _02826_ VGND VGND VPWR VPWR _02827_ sky130_fd_sc_hd__clkbuf_4
X_18116_ net179 _02396_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18047_ net1220 _02327_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_15259_ _05441_ VGND VGND VPWR VPWR _02758_ sky130_fd_sc_hd__buf_4
XFILLER_0_100_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09820_ _05481_ VGND VGND VPWR VPWR _02515_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09751_ _05439_ VGND VGND VPWR VPWR _05440_ sky130_fd_sc_hd__clkbuf_4
X_08702_ _04421_ _04420_ _04282_ VGND VGND VPWR VPWR _04422_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_107_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09682_ _05371_ _05372_ _05373_ _04708_ VGND VGND VPWR VPWR _05374_ sky130_fd_sc_hd__o31a_1
XFILLER_0_146_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08633_ _04234_ _04352_ VGND VGND VPWR VPWR _04353_ sky130_fd_sc_hd__and2_1
XFILLER_0_55_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08564_ CPU.mem_wdata\[4\] CPU.Iimm\[4\] _04203_ VGND VGND VPWR VPWR _04284_ sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_120_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08495_ CPU.Jimm\[13\] VGND VGND VPWR VPWR _04215_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09116_ CPU.PC\[20\] _04826_ VGND VGND VPWR VPWR _04828_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_135_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09047_ _04761_ VGND VGND VPWR VPWR _04762_ sky130_fd_sc_hd__buf_4
XFILLER_0_20_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold450 CPU.PC\[19\] VGND VGND VPWR VPWR net1691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 CPU.registerFile\[14\]\[24\] VGND VGND VPWR VPWR net1702 sky130_fd_sc_hd__dlygate4sd3_1
X_14960__1038 clknet_1_1__leaf__02711_ VGND VGND VPWR VPWR net1070 sky130_fd_sc_hd__inv_2
Xhold472 per_uart.uart0.txd_reg\[1\] VGND VGND VPWR VPWR net1713 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold483 CPU.registerFile\[1\]\[5\] VGND VGND VPWR VPWR net1724 sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 CPU.registerFile\[19\]\[29\] VGND VGND VPWR VPWR net1735 sky130_fd_sc_hd__dlygate4sd3_1
X_15182__1207 clknet_1_0__leaf__02748_ VGND VGND VPWR VPWR net1239 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_5_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09949_ _05566_ VGND VGND VPWR VPWR _02471_ sky130_fd_sc_hd__clkbuf_1
X_12960_ _07398_ _07400_ VGND VGND VPWR VPWR _07401_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_51_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1150 CPU.registerFile\[9\]\[29\] VGND VGND VPWR VPWR net2391 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11911_ _06721_ VGND VGND VPWR VPWR _01614_ sky130_fd_sc_hd__clkbuf_1
Xhold1161 CPU.registerFile\[25\]\[31\] VGND VGND VPWR VPWR net2402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1172 CPU.registerFile\[23\]\[11\] VGND VGND VPWR VPWR net2413 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1183 CPU.registerFile\[11\]\[28\] VGND VGND VPWR VPWR net2424 sky130_fd_sc_hd__dlygate4sd3_1
X_12891_ _07324_ _07328_ _07329_ _07332_ VGND VGND VPWR VPWR _07333_ sky130_fd_sc_hd__a22o_1
Xhold1194 CPU.aluReg\[3\] VGND VGND VPWR VPWR net2435 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_301 _07333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14543__662 clknet_1_0__leaf__02670_ VGND VGND VPWR VPWR net694 sky130_fd_sc_hd__inv_2
XANTENNA_312 _07914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11842_ net2091 _05689_ _06675_ VGND VGND VPWR VPWR _06685_ sky130_fd_sc_hd__mux2_1
XANTENNA_323 _07914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_334 _02861_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_345 _05338_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_356 _07268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_367 _02889_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11773_ _06648_ VGND VGND VPWR VPWR _01679_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_378 _07318_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_389 _07271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_16300_ CPU.registerFile\[1\]\[26\] _02867_ _03772_ _02895_ VGND VGND VPWR VPWR _03773_
+ sky130_fd_sc_hd__a22o_1
X_13512_ _07380_ _07932_ _07936_ _07646_ VGND VGND VPWR VPWR _07937_ sky130_fd_sc_hd__o211a_1
X_17280_ net469 _01568_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_10724_ _06055_ VGND VGND VPWR VPWR _02138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_155_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16231_ _03701_ _03705_ _08410_ VGND VGND VPWR VPWR _03706_ sky130_fd_sc_hd__a21o_1
X_13443_ _07866_ _07869_ _07584_ VGND VGND VPWR VPWR _07870_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_137_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10655_ _05965_ _05962_ net2 VGND VGND VPWR VPWR _00004_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_153_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14199__377 clknet_1_0__leaf__08429_ VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__inv_2
XFILLER_0_23_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16162_ _02914_ _03638_ _02965_ VGND VGND VPWR VPWR _03639_ sky130_fd_sc_hd__a21o_1
X_13374_ CPU.registerFile\[2\]\[14\] _07322_ VGND VGND VPWR VPWR _07803_ sky130_fd_sc_hd__or2_1
Xclkload17 clknet_leaf_23_clk VGND VGND VPWR VPWR clkload17/Y sky130_fd_sc_hd__clkinv_1
Xclkload28 clknet_1_0__leaf__02749_ VGND VGND VPWR VPWR clkload28/X sky130_fd_sc_hd__clkbuf_8
X_10586_ net1476 _05968_ _05974_ _05936_ VGND VGND VPWR VPWR _02194_ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload39 clknet_1_0__leaf__02746_ VGND VGND VPWR VPWR clkload39/Y sky130_fd_sc_hd__clkinvlp_4
X_12325_ _04696_ net2119 _06977_ VGND VGND VPWR VPWR _06979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16093_ CPU.registerFile\[22\]\[20\] _08399_ VGND VGND VPWR VPWR _03572_ sky130_fd_sc_hd__and2_1
XFILLER_0_121_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12256_ _06859_ VGND VGND VPWR VPWR _06927_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_71_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11207_ _06312_ VGND VGND VPWR VPWR _01912_ sky130_fd_sc_hd__clkbuf_1
X_12187_ CPU.aluReg\[30\] _06871_ _06873_ VGND VGND VPWR VPWR _06874_ sky130_fd_sc_hd__a21o_1
X_11138_ CPU.registerFile\[8\]\[10\] _05715_ _06274_ VGND VGND VPWR VPWR _06276_ sky130_fd_sc_hd__mux2_1
X_16995_ clknet_leaf_28_clk _01321_ VGND VGND VPWR VPWR CPU.rs2\[26\] sky130_fd_sc_hd__dfxtp_1
X_14626__737 clknet_1_1__leaf__02678_ VGND VGND VPWR VPWR net769 sky130_fd_sc_hd__inv_2
X_11069_ net2506 _05715_ _06237_ VGND VGND VPWR VPWR _06239_ sky130_fd_sc_hd__mux2_1
X_15946_ _08411_ _03421_ _03429_ _02993_ VGND VGND VPWR VPWR _03430_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_0_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_8
X_15877_ _02948_ _03359_ _03362_ VGND VGND VPWR VPWR _03363_ sky130_fd_sc_hd__or3_2
XFILLER_0_116_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17616_ net805 _01904_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_552 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17547_ net736 _01835_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_451 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17478_ net667 _01766_ VGND VGND VPWR VPWR mapped_spi_flash.div_counter\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16429_ CPU.registerFile\[9\]\[30\] CPU.registerFile\[13\]\[30\] _02798_ VGND VGND
+ VPWR VPWR _03898_ sky130_fd_sc_hd__mux2_1
X_14672__779 clknet_1_1__leaf__02682_ VGND VGND VPWR VPWR net811 sky130_fd_sc_hd__inv_2
XFILLER_0_42_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16541__17 clknet_1_1__leaf__03965_ VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__inv_2
XFILLER_0_124_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_113_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09803_ _05472_ VGND VGND VPWR VPWR _02523_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09734_ _05420_ _05423_ _04708_ VGND VGND VPWR VPWR _05424_ sky130_fd_sc_hd__o21a_1
X_09665_ CPU.cycles\[4\] _04687_ _05342_ _05357_ VGND VGND VPWR VPWR _05358_ sky130_fd_sc_hd__a211o_2
XFILLER_0_97_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08616_ _04335_ _04253_ VGND VGND VPWR VPWR _04336_ sky130_fd_sc_hd__nand2_2
X_09596_ CPU.PC\[6\] VGND VGND VPWR VPWR _05291_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08547_ _04266_ VGND VGND VPWR VPWR _04267_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08478_ CPU.instr\[2\] net1275 VGND VGND VPWR VPWR _04198_ sky130_fd_sc_hd__or2b_4
XFILLER_0_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10440_ net1374 _05849_ _05858_ _05855_ VGND VGND VPWR VPWR _02224_ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_150_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10371_ _05807_ VGND VGND VPWR VPWR _02243_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12110_ _04798_ net2005 _06819_ VGND VGND VPWR VPWR _06827_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13090_ CPU.registerFile\[28\]\[5\] CPU.registerFile\[24\]\[5\] _07352_ VGND VGND
+ VPWR VPWR _07528_ sky130_fd_sc_hd__mux2_1
X_12041_ _06790_ VGND VGND VPWR VPWR _01552_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_53_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold280 mapped_spi_ram.snd_bitcount\[1\] VGND VGND VPWR VPWR net1521 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold291 CPU.rs2\[12\] VGND VGND VPWR VPWR net1532 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15800_ CPU.registerFile\[1\]\[11\] _02814_ _03287_ _02943_ VGND VGND VPWR VPWR _03288_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_148_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16780_ _04052_ _05005_ _08453_ VGND VGND VPWR VPWR _04093_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_29_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12943_ CPU.registerFile\[16\]\[2\] CPU.registerFile\[20\]\[2\] _07339_ VGND VGND
+ VPWR VPWR _07384_ sky130_fd_sc_hd__mux2_1
X_15731_ CPU.registerFile\[16\]\[9\] CPU.registerFile\[18\]\[9\] _03032_ VGND VGND
+ VPWR VPWR _03221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12874_ _07312_ _07313_ _07315_ VGND VGND VPWR VPWR _07316_ sky130_fd_sc_hd__mux2_1
XANTENNA_120 _05524_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15662_ CPU.registerFile\[18\]\[7\] _02832_ _02835_ CPU.registerFile\[19\]\[7\] _03074_
+ VGND VGND VPWR VPWR _03154_ sky130_fd_sc_hd__o221a_1
XFILLER_0_158_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_131 _05549_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_142 _05719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17401_ net590 _01689_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_bitcount\[1\] sky130_fd_sc_hd__dfxtp_1
X_11825_ _06676_ VGND VGND VPWR VPWR _01655_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_153 _07271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15593_ _02759_ _03083_ _03085_ _02767_ VGND VGND VPWR VPWR _03086_ sky130_fd_sc_hd__a211o_1
XANTENNA_164 _07322_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_175 _07476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_186 _07799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_197 _07841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17332_ net521 _01620_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_11756_ _04659_ net1769 _06639_ VGND VGND VPWR VPWR _06640_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__03970_ clknet_0__03970_ VGND VGND VPWR VPWR clknet_1_1__leaf__03970_
+ sky130_fd_sc_hd__clkbuf_16
X_14207__384 clknet_1_0__leaf__08430_ VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__inv_2
XFILLER_0_138_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14814__907 clknet_1_1__leaf__02696_ VGND VGND VPWR VPWR net939 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_64_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10707_ _05514_ net1661 _06045_ VGND VGND VPWR VPWR _06047_ sky130_fd_sc_hd__mux2_1
X_17263_ net453 _01551_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11687_ net1424 _06590_ _06596_ _06594_ VGND VGND VPWR VPWR _01712_ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_125_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13426_ _07519_ _07852_ _07853_ VGND VGND VPWR VPWR _07854_ sky130_fd_sc_hd__o21a_1
X_16214_ CPU.registerFile\[27\]\[23\] CPU.registerFile\[31\]\[23\] _02798_ VGND VGND
+ VPWR VPWR _03690_ sky130_fd_sc_hd__mux2_1
X_17194_ clknet_leaf_25_clk _01482_ VGND VGND VPWR VPWR CPU.Iimm\[4\] sky130_fd_sc_hd__dfxtp_1
X_10638_ net1486 _05996_ _06003_ _05993_ VGND VGND VPWR VPWR _02171_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload106 clknet_1_0__leaf__08359_ VGND VGND VPWR VPWR clkload106/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_153_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12754__207 clknet_1_0__leaf__07221_ VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__inv_2
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload117 clknet_1_0__leaf__03965_ VGND VGND VPWR VPWR clkload117/Y sky130_fd_sc_hd__clkinvlp_4
X_16145_ CPU.registerFile\[20\]\[21\] CPU.registerFile\[21\]\[21\] _08394_ VGND VGND
+ VPWR VPWR _03623_ sky130_fd_sc_hd__mux2_1
X_13357_ CPU.registerFile\[23\]\[13\] _07276_ _07277_ CPU.registerFile\[19\]\[13\]
+ _07278_ VGND VGND VPWR VPWR _07787_ sky130_fd_sc_hd__o221a_1
X_10569_ _05961_ VGND VGND VPWR VPWR _02198_ sky130_fd_sc_hd__clkbuf_1
X_13999__280 clknet_1_0__leaf__08360_ VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__inv_2
XFILLER_0_87_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12308_ _06966_ VGND VGND VPWR VPWR _01427_ sky130_fd_sc_hd__clkbuf_1
X_16076_ CPU.registerFile\[31\]\[19\] _03072_ VGND VGND VPWR VPWR _03556_ sky130_fd_sc_hd__or2_1
X_13288_ _07360_ _07716_ _07719_ _07392_ VGND VGND VPWR VPWR _07720_ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12239_ CPU.aluIn1\[19\] _06913_ _06894_ VGND VGND VPWR VPWR _06914_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16978_ clknet_leaf_26_clk _01304_ VGND VGND VPWR VPWR CPU.rs2\[9\] sky130_fd_sc_hd__dfxtp_1
Xinput4 spi_miso_ram VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
X_15929_ _03406_ _03412_ _02879_ VGND VGND VPWR VPWR _03413_ sky130_fd_sc_hd__o21a_1
XFILLER_0_127_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09450_ _05151_ VGND VGND VPWR VPWR _02563_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_2_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_84_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09381_ CPU.PC\[15\] _04924_ CPU.PC\[16\] VGND VGND VPWR VPWR _05086_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15181__1206 clknet_1_0__leaf__02748_ VGND VGND VPWR VPWR net1238 sky130_fd_sc_hd__inv_2
XFILLER_0_7_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_132_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15196__109 clknet_1_0__leaf__02750_ VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__inv_2
XFILLER_0_77_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14609__721 clknet_1_0__leaf__02677_ VGND VGND VPWR VPWR net753 sky130_fd_sc_hd__inv_2
X_09717_ mapped_spi_ram.rcv_data\[25\] net17 _04643_ per_uart.rx_data\[1\] _05277_
+ VGND VGND VPWR VPWR _05407_ sky130_fd_sc_hd__a221o_1
X_09648_ _05338_ _05281_ _05340_ _05277_ VGND VGND VPWR VPWR _05341_ sky130_fd_sc_hd__o22a_1
XFILLER_0_69_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_139_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09579_ _05274_ VGND VGND VPWR VPWR _02557_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11610_ net1373 _06501_ _06496_ CPU.mem_wdata\[3\] _06508_ VGND VGND VPWR VPWR _06544_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12590_ _07118_ VGND VGND VPWR VPWR _01264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11541_ CPU.mem_rstrb _04783_ _06493_ VGND VGND VPWR VPWR _06496_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_25_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14655__763 clknet_1_0__leaf__02681_ VGND VGND VPWR VPWR net795 sky130_fd_sc_hd__inv_2
XFILLER_0_34_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14260_ _05247_ _05261_ _05297_ _08438_ VGND VGND VPWR VPWR _08439_ sky130_fd_sc_hd__or4_1
X_11472_ _05528_ net2430 _06444_ VGND VGND VPWR VPWR _06453_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13211_ _07639_ _07642_ _07643_ _07644_ _07570_ VGND VGND VPWR VPWR _07645_ sky130_fd_sc_hd__a221o_1
XFILLER_0_107_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10423_ net2425 _05825_ _05827_ mapped_spi_flash.cmd_addr\[23\] VGND VGND VPWR VPWR
+ _05845_ sky130_fd_sc_hd__a22o_1
X_14191_ clknet_1_0__leaf__08363_ VGND VGND VPWR VPWR _08429_ sky130_fd_sc_hd__buf_1
X_13142_ CPU.registerFile\[5\]\[7\] CPU.registerFile\[4\]\[7\] _07577_ VGND VGND VPWR
+ VPWR _07578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10354_ _05798_ VGND VGND VPWR VPWR _02251_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13073_ CPU.registerFile\[5\]\[5\] CPU.registerFile\[4\]\[5\] net14 VGND VGND VPWR
+ VPWR _07511_ sky130_fd_sc_hd__mux2_1
X_17950_ net1139 _02234_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[30\] sky130_fd_sc_hd__dfxtp_1
X_10285_ _05761_ VGND VGND VPWR VPWR _02298_ sky130_fd_sc_hd__clkbuf_1
X_14053__329 clknet_1_1__leaf__08365_ VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__inv_2
X_12024_ _05448_ net2049 _06746_ VGND VGND VPWR VPWR _06781_ sky130_fd_sc_hd__mux2_1
X_16901_ net1536 _04177_ VGND VGND VPWR VPWR _04178_ sky130_fd_sc_hd__or2_1
X_17881_ net1070 net1338 VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dfxtp_1
X_16832_ per_uart.uart0.tx_bitcount\[1\] per_uart.uart0.tx_bitcount\[0\] per_uart.uart0.tx_bitcount\[2\]
+ VGND VGND VPWR VPWR _04132_ sky130_fd_sc_hd__a21oi_1
X_14820__911 clknet_1_0__leaf__02698_ VGND VGND VPWR VPWR net943 sky130_fd_sc_hd__inv_2
X_16763_ _04001_ _05055_ _03990_ VGND VGND VPWR VPWR _04079_ sky130_fd_sc_hd__a21o_1
X_15714_ CPU.registerFile\[2\]\[9\] _02872_ _02873_ CPU.registerFile\[3\]\[9\] _02875_
+ VGND VGND VPWR VPWR _03204_ sky130_fd_sc_hd__a221o_1
X_12926_ CPU.registerFile\[23\]\[2\] _07362_ _07363_ CPU.registerFile\[19\]\[2\] _07366_
+ VGND VGND VPWR VPWR _07367_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_66_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16694_ _04016_ _04020_ _05942_ VGND VGND VPWR VPWR _02586_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_66_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15645_ _02797_ _03134_ _03135_ _03136_ _03054_ VGND VGND VPWR VPWR _03137_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12857_ _04971_ VGND VGND VPWR VPWR _07300_ sky130_fd_sc_hd__buf_4
XFILLER_0_158_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14738__838 clknet_1_0__leaf__02689_ VGND VGND VPWR VPWR net870 sky130_fd_sc_hd__inv_2
XFILLER_0_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11808_ _05306_ net2530 _06661_ VGND VGND VPWR VPWR _06667_ sky130_fd_sc_hd__mux2_1
X_18364_ clknet_leaf_3_clk _02642_ VGND VGND VPWR VPWR per_uart.d_in_uart\[4\] sky130_fd_sc_hd__dfxtp_1
X_12788_ _05232_ VGND VGND VPWR VPWR _07231_ sky130_fd_sc_hd__clkbuf_4
X_15576_ CPU.registerFile\[16\]\[5\] _03068_ _03069_ CPU.registerFile\[17\]\[5\] _02779_
+ VGND VGND VPWR VPWR _03070_ sky130_fd_sc_hd__o221a_1
XFILLER_0_17_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17315_ net504 _01603_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_11739_ _06628_ VGND VGND VPWR VPWR _01693_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18295_ net128 _02575_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17246_ net436 _01534_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13409_ CPU.registerFile\[23\]\[15\] _07629_ _07488_ CPU.registerFile\[19\]\[15\]
+ _07836_ VGND VGND VPWR VPWR _07837_ sky130_fd_sc_hd__o221a_1
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17177_ clknet_leaf_25_clk _01465_ VGND VGND VPWR VPWR CPU.Bimm\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16128_ _02797_ _03603_ _03604_ _03605_ _02807_ VGND VGND VPWR VPWR _03606_ sky130_fd_sc_hd__a221o_1
XFILLER_0_141_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08950_ _04669_ VGND VGND VPWR VPWR _02581_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_94_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16059_ CPU.registerFile\[20\]\[19\] _02855_ _03026_ VGND VGND VPWR VPWR _03539_
+ sky130_fd_sc_hd__a21o_1
Xclkbuf_1_1__f__02697_ clknet_0__02697_ VGND VGND VPWR VPWR clknet_1_1__leaf__02697_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_110_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__07224_ clknet_0__07224_ VGND VGND VPWR VPWR clknet_1_1__leaf__07224_
+ sky130_fd_sc_hd__clkbuf_16
X_08881_ CPU.PC\[16\] _04598_ _04600_ _04562_ VGND VGND VPWR VPWR _04601_ sky130_fd_sc_hd__a22oi_4
XPHY_EDGE_ROW_135_Right_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09502_ _04430_ _05200_ VGND VGND VPWR VPWR _05201_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09433_ _04216_ _05132_ _05133_ _05134_ _04717_ VGND VGND VPWR VPWR _05135_ sky130_fd_sc_hd__o221a_1
XFILLER_0_94_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09364_ mapped_spi_ram.rcv_data\[8\] net16 _04690_ mapped_spi_flash.rcv_data\[8\]
+ VGND VGND VPWR VPWR _05069_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_20 _02926_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_09295_ CPU.PC\[20\] _04927_ VGND VGND VPWR VPWR _05004_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_31 _03072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_42 _03941_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_53 _04958_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_64 _05065_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_75 _05169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_86 _05284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_97 _05359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15204__116 clknet_1_0__leaf__02751_ VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__inv_2
XFILLER_0_100_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10070_ _05630_ VGND VGND VPWR VPWR _02382_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_102_Right_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_145_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__08431_ clknet_0__08431_ VGND VGND VPWR VPWR clknet_1_0__leaf__08431_
+ sky130_fd_sc_hd__clkbuf_16
Xmax_cap22 net23 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
X_13760_ CPU.registerFile\[6\]\[26\] CPU.registerFile\[7\]\[26\] _07641_ VGND VGND
+ VPWR VPWR _08177_ sky130_fd_sc_hd__mux2_1
X_10972_ _06187_ VGND VGND VPWR VPWR _02022_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_39_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__08362_ clknet_0__08362_ VGND VGND VPWR VPWR clknet_1_0__leaf__08362_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_39_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12711_ per_uart.uart0.enable16_counter\[14\] _07192_ VGND VGND VPWR VPWR _07193_
+ sky130_fd_sc_hd__or2_1
X_13691_ _07584_ _08103_ _08110_ _07703_ VGND VGND VPWR VPWR _08111_ sky130_fd_sc_hd__a31o_1
XFILLER_0_97_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15250__158 clknet_1_0__leaf__02755_ VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__inv_2
XFILLER_0_155_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12642_ net1439 _07144_ VGND VGND VPWR VPWR _07147_ sky130_fd_sc_hd__nor2_1
X_15430_ CPU.registerFile\[29\]\[2\] _02926_ VGND VGND VPWR VPWR _02927_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15361_ CPU.registerFile\[14\]\[1\] CPU.registerFile\[10\]\[1\] _02761_ VGND VGND
+ VPWR VPWR _02859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12573_ CPU.registerFile\[4\]\[9\] _05229_ _07107_ VGND VGND VPWR VPWR _07110_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17100_ net358 _01422_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11524_ _06483_ net21 mapped_spi_ram.state\[1\] VGND VGND VPWR VPWR _06486_ sky130_fd_sc_hd__o21a_1
X_15292_ _02772_ VGND VGND VPWR VPWR _02791_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_124_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18080_ net143 _02360_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17031_ net289 _01353_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_11455_ _06432_ VGND VGND VPWR VPWR _06444_ sky130_fd_sc_hd__buf_4
XFILLER_0_135_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_12_Left_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__02720_ _02720_ VGND VGND VPWR VPWR clknet_0__02720_ sky130_fd_sc_hd__clkbuf_16
X_10406_ _05830_ _05833_ VGND VGND VPWR VPWR _05834_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14174_ _08424_ VGND VGND VPWR VPWR _01487_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11386_ _06407_ VGND VGND VPWR VPWR _01828_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13125_ CPU.registerFile\[30\]\[6\] CPU.registerFile\[26\]\[6\] _07352_ VGND VGND
+ VPWR VPWR _07562_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10337_ _05514_ net2302 _05788_ VGND VGND VPWR VPWR _05790_ sky130_fd_sc_hd__mux2_1
X_13056_ _07475_ _07493_ _07494_ VGND VGND VPWR VPWR _07495_ sky130_fd_sc_hd__o21a_1
X_17933_ net1122 _02217_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[13\] sky130_fd_sc_hd__dfxtp_1
X_10268_ _05514_ net2459 _05751_ VGND VGND VPWR VPWR _05753_ sky130_fd_sc_hd__mux2_1
X_15180__1205 clknet_1_0__leaf__02748_ VGND VGND VPWR VPWR net1237 sky130_fd_sc_hd__inv_2
X_12007_ _06772_ VGND VGND VPWR VPWR _01569_ sky130_fd_sc_hd__clkbuf_1
X_17864_ net1053 _02148_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_10199_ CPU.registerFile\[1\]\[13\] _05708_ _05692_ VGND VGND VPWR VPWR _05709_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16815_ _05830_ _04119_ VGND VGND VPWR VPWR _04120_ sky130_fd_sc_hd__and2_1
X_17795_ net984 _02079_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[17\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_21_Left_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16746_ _04050_ _04062_ _04063_ _04064_ VGND VGND VPWR VPWR _04065_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_17_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12909_ _07291_ VGND VGND VPWR VPWR _07351_ sky130_fd_sc_hd__clkbuf_4
X_14326__467 clknet_1_1__leaf__08465_ VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__inv_2
XFILLER_0_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16677_ _08453_ VGND VGND VPWR VPWR _04006_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_88_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13889_ _08297_ _08298_ _08299_ _08301_ VGND VGND VPWR VPWR _08302_ sky130_fd_sc_hd__a22o_2
XFILLER_0_75_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15628_ CPU.registerFile\[8\]\[7\] _02763_ _03117_ _03119_ VGND VGND VPWR VPWR _03120_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13964__249 clknet_1_1__leaf__08356_ VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__inv_2
XFILLER_0_72_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18347_ clknet_leaf_1_clk _02627_ VGND VGND VPWR VPWR per_uart.uart0.rx_count16\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15559_ CPU.registerFile\[25\]\[5\] _02802_ _02803_ VGND VGND VPWR VPWR _03053_ sky130_fd_sc_hd__o21a_1
X_09080_ CPU.aluIn1\[24\] _04235_ _04209_ VGND VGND VPWR VPWR _04793_ sky130_fd_sc_hd__o21a_1
XFILLER_0_72_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18278_ net111 _02558_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17229_ net419 _01517_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_96_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__03967_ _03967_ VGND VGND VPWR VPWR clknet_0__03967_ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_96_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold802 CPU.registerFile\[29\]\[14\] VGND VGND VPWR VPWR net2043 sky130_fd_sc_hd__dlygate4sd3_1
Xhold813 CPU.registerFile\[3\]\[17\] VGND VGND VPWR VPWR net2054 sky130_fd_sc_hd__dlygate4sd3_1
Xhold824 CPU.registerFile\[12\]\[10\] VGND VGND VPWR VPWR net2065 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold835 CPU.registerFile\[27\]\[20\] VGND VGND VPWR VPWR net2076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 CPU.registerFile\[13\]\[23\] VGND VGND VPWR VPWR net2087 sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 CPU.registerFile\[6\]\[26\] VGND VGND VPWR VPWR net2098 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold868 per_uart.uart0.rx_bitcount\[1\] VGND VGND VPWR VPWR net2109 sky130_fd_sc_hd__dlygate4sd3_1
X_09982_ _05537_ net2186 _05581_ VGND VGND VPWR VPWR _05584_ sky130_fd_sc_hd__mux2_1
Xhold879 CPU.registerFile\[13\]\[4\] VGND VGND VPWR VPWR net2120 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__02749_ clknet_0__02749_ VGND VGND VPWR VPWR clknet_1_1__leaf__02749_
+ sky130_fd_sc_hd__clkbuf_16
X_14036__313 clknet_1_1__leaf__08364_ VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__inv_2
Xclkbuf_0__08356_ _08356_ VGND VGND VPWR VPWR clknet_0__08356_ sky130_fd_sc_hd__clkbuf_16
X_08933_ _04499_ CPU.instr\[2\] _04291_ VGND VGND VPWR VPWR _04653_ sky130_fd_sc_hd__or3_1
XFILLER_0_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12767__217 clknet_1_1__leaf__07224_ VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__inv_2
X_08864_ _04577_ _04583_ _04579_ VGND VGND VPWR VPWR _04584_ sky130_fd_sc_hd__and3_1
XFILLER_0_99_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08795_ _04513_ _04514_ VGND VGND VPWR VPWR _04515_ sky130_fd_sc_hd__nor2_1
X_16646__90 clknet_1_0__leaf__03989_ VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_140_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_820 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09416_ _04437_ _04396_ _04436_ VGND VGND VPWR VPWR _05119_ sky130_fd_sc_hd__or3_1
XFILLER_0_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14082__355 clknet_1_1__leaf__08368_ VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__inv_2
XFILLER_0_48_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09347_ _04442_ _04390_ _04441_ VGND VGND VPWR VPWR _05053_ sky130_fd_sc_hd__or3_1
XFILLER_0_47_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09278_ _04986_ VGND VGND VPWR VPWR _04987_ sky130_fd_sc_hd__buf_4
XFILLER_0_106_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11240_ net1628 _05681_ _06324_ VGND VGND VPWR VPWR _06330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11171_ _06293_ VGND VGND VPWR VPWR _01929_ sky130_fd_sc_hd__clkbuf_1
X_14767__864 clknet_1_0__leaf__02692_ VGND VGND VPWR VPWR net896 sky130_fd_sc_hd__inv_2
X_10122_ net2038 _05253_ _05655_ VGND VGND VPWR VPWR _05659_ sky130_fd_sc_hd__mux2_1
X_16527__194 clknet_1_1__leaf__03964_ VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__inv_2
X_10053_ net2463 _05253_ _05618_ VGND VGND VPWR VPWR _05622_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13812_ CPU.registerFile\[31\]\[27\] _07556_ _07557_ CPU.registerFile\[27\]\[27\]
+ _08227_ VGND VGND VPWR VPWR _08228_ sky130_fd_sc_hd__o221a_1
X_17580_ net769 _01868_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[30\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_3_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10955_ _05631_ _06141_ VGND VGND VPWR VPWR _06178_ sky130_fd_sc_hd__nor2_4
X_13743_ CPU.registerFile\[19\]\[25\] _07619_ _08160_ VGND VGND VPWR VPWR _08161_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16462_ CPU.registerFile\[6\]\[31\] _02828_ VGND VGND VPWR VPWR _03930_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13674_ CPU.registerFile\[19\]\[23\] _07383_ _08093_ _07254_ VGND VGND VPWR VPWR
+ _08094_ sky130_fd_sc_hd__o211a_1
X_10886_ _04665_ _04663_ _04664_ CPU.writeBack VGND VGND VPWR VPWR _06141_ sky130_fd_sc_hd__or4bb_4
XTAP_TAPCELL_ROW_158_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18201_ net42 _02481_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_158_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15413_ _05441_ VGND VGND VPWR VPWR _02910_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_158_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_503 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12625_ CPU.cycles\[0\] CPU.cycles\[1\] net1419 VGND VGND VPWR VPWR _07137_ sky130_fd_sc_hd__a21oi_1
X_16393_ CPU.registerFile\[5\]\[29\] CPU.registerFile\[4\]\[29\] _05092_ VGND VGND
+ VPWR VPWR _03863_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18132_ net195 _02412_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_12556_ CPU.registerFile\[4\]\[17\] _05065_ _07096_ VGND VGND VPWR VPWR _07101_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15344_ _05029_ VGND VGND VPWR VPWR _02843_ sky130_fd_sc_hd__buf_4
XFILLER_0_81_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11507_ mapped_spi_ram.state\[2\] CPU.mem_rstrb _05068_ VGND VGND VPWR VPWR _06474_
+ sky130_fd_sc_hd__and3_2
X_18063_ net1236 _02343_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12487_ _07064_ VGND VGND VPWR VPWR _01346_ sky130_fd_sc_hd__clkbuf_1
X_15275_ CPU.registerFile\[15\]\[0\] CPU.registerFile\[11\]\[0\] _02773_ VGND VGND
+ VPWR VPWR _02774_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17014_ net272 _01336_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold109 mapped_spi_ram.cmd_addr\[7\] VGND VGND VPWR VPWR net1350 sky130_fd_sc_hd__dlygate4sd3_1
X_11438_ _06435_ VGND VGND VPWR VPWR _01804_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__02703_ _02703_ VGND VGND VPWR VPWR clknet_0__02703_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14157_ _08415_ VGND VGND VPWR VPWR _01479_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11369_ _05493_ net1856 _06397_ VGND VGND VPWR VPWR _06399_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_74_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13108_ _04939_ _07542_ _07544_ _04972_ VGND VGND VPWR VPWR _07545_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_91_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14088_ _07128_ _08369_ _05275_ _05112_ VGND VGND VPWR VPWR _08370_ sky130_fd_sc_hd__and4b_1
X_13039_ CPU.registerFile\[29\]\[4\] _07325_ _07326_ CPU.registerFile\[25\]\[4\] _07249_
+ VGND VGND VPWR VPWR _07478_ sky130_fd_sc_hd__o221a_1
XFILLER_0_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17916_ net1105 _02200_ VGND VGND VPWR VPWR mapped_spi_flash.snd_bitcount\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17847_ net1036 _02131_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_08580_ _04290_ _04297_ _04299_ VGND VGND VPWR VPWR _04300_ sky130_fd_sc_hd__nand3_2
X_17778_ net967 _02062_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_15162__1189 clknet_1_1__leaf__02746_ VGND VGND VPWR VPWR net1221 sky130_fd_sc_hd__inv_2
X_16729_ _05289_ VGND VGND VPWR VPWR _04050_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_105_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15233__142 clknet_1_1__leaf__02754_ VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_122_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09201_ _04910_ _04912_ VGND VGND VPWR VPWR _04913_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09132_ CPU.Jimm\[15\] _04829_ _04831_ VGND VGND VPWR VPWR _04844_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09063_ _04655_ VGND VGND VPWR VPWR _04777_ sky130_fd_sc_hd__buf_6
XFILLER_0_142_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold610 CPU.registerFile\[30\]\[29\] VGND VGND VPWR VPWR net1851 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold621 CPU.registerFile\[10\]\[27\] VGND VGND VPWR VPWR net1862 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold632 CPU.registerFile\[22\]\[0\] VGND VGND VPWR VPWR net1873 sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 CPU.registerFile\[12\]\[17\] VGND VGND VPWR VPWR net1884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold654 CPU.registerFile\[4\]\[21\] VGND VGND VPWR VPWR net1895 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold665 CPU.registerFile\[27\]\[5\] VGND VGND VPWR VPWR net1906 sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 CPU.registerFile\[25\]\[4\] VGND VGND VPWR VPWR net1917 sky130_fd_sc_hd__dlygate4sd3_1
Xhold687 CPU.registerFile\[13\]\[21\] VGND VGND VPWR VPWR net1928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold698 CPU.registerFile\[16\]\[15\] VGND VGND VPWR VPWR net1939 sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ _05520_ net1784 _05570_ VGND VGND VPWR VPWR _05575_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08916_ _04621_ VGND VGND VPWR VPWR _04636_ sky130_fd_sc_hd__inv_2
X_09896_ _05187_ VGND VGND VPWR VPWR _05532_ sky130_fd_sc_hd__buf_4
XFILLER_0_99_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08847_ CPU.aluIn1\[18\] _04494_ VGND VGND VPWR VPWR _04567_ sky130_fd_sc_hd__or2_1
X_08778_ _04497_ VGND VGND VPWR VPWR _04498_ sky130_fd_sc_hd__buf_2
X_14309__451 clknet_1_0__leaf__08464_ VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10740_ _05547_ net2337 _06056_ VGND VGND VPWR VPWR _06064_ sky130_fd_sc_hd__mux2_1
X_13947__233 clknet_1_0__leaf__07226_ VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__inv_2
XFILLER_0_137_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10671_ mapped_spi_flash.rcv_bitcount\[1\] mapped_spi_flash.rcv_bitcount\[0\] net1357
+ VGND VGND VPWR VPWR _06026_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_138_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12410_ _07023_ VGND VGND VPWR VPWR _01382_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13390_ CPU.registerFile\[14\]\[14\] CPU.registerFile\[10\]\[14\] _07274_ VGND VGND
+ VPWR VPWR _07819_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14008__289 clknet_1_1__leaf__08360_ VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__inv_2
XFILLER_0_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12341_ _04958_ net1811 _06977_ VGND VGND VPWR VPWR _06987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14201__379 clknet_1_0__leaf__08429_ VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__inv_2
X_12272_ _06870_ VGND VGND VPWR VPWR _06939_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11223_ _06320_ VGND VGND VPWR VPWR _01904_ sky130_fd_sc_hd__clkbuf_1
X_14355__493 clknet_1_1__leaf__08468_ VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__inv_2
XFILLER_0_31_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11154_ net2488 _05731_ _06274_ VGND VGND VPWR VPWR _06284_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13993__275 clknet_1_1__leaf__08359_ VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__inv_2
X_10105_ net2383 _05090_ _05644_ VGND VGND VPWR VPWR _05650_ sky130_fd_sc_hd__mux2_1
X_11085_ net1979 _05731_ _06237_ VGND VGND VPWR VPWR _06247_ sky130_fd_sc_hd__mux2_1
X_15962_ CPU.registerFile\[29\]\[16\] _02918_ VGND VGND VPWR VPWR _03445_ sky130_fd_sc_hd__or2_1
X_17701_ net890 _01989_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_10036_ net2037 _05090_ _05607_ VGND VGND VPWR VPWR _05613_ sky130_fd_sc_hd__mux2_1
X_15893_ _02911_ _03375_ _03377_ _02794_ VGND VGND VPWR VPWR _03378_ sky130_fd_sc_hd__a211o_1
X_17632_ net821 _01920_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_904 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16625__71 clknet_1_1__leaf__03971_ VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__inv_2
X_17563_ net752 _01851_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_11987_ _05046_ net1682 _06758_ VGND VGND VPWR VPWR _06762_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13726_ _07305_ _08143_ VGND VGND VPWR VPWR _08144_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_27_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10938_ _06169_ VGND VGND VPWR VPWR _02038_ sky130_fd_sc_hd__clkbuf_1
X_17494_ net683 _01782_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14520__641 clknet_1_1__leaf__02668_ VGND VGND VPWR VPWR net673 sky130_fd_sc_hd__inv_2
X_16640__85 clknet_1_0__leaf__03988_ VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_27_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16445_ _03912_ _03913_ _08400_ VGND VGND VPWR VPWR _03914_ sky130_fd_sc_hd__mux2_1
X_10869_ _06132_ VGND VGND VPWR VPWR _02070_ sky130_fd_sc_hd__clkbuf_1
X_13657_ _07334_ _08067_ _08070_ _08077_ _07766_ VGND VGND VPWR VPWR _08078_ sky130_fd_sc_hd__o311a_1
XFILLER_0_38_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12608_ _04589_ _07126_ VGND VGND VPWR VPWR _07127_ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16376_ _03842_ _03846_ _02949_ VGND VGND VPWR VPWR _03847_ sky130_fd_sc_hd__a21o_1
X_13588_ CPU.registerFile\[28\]\[20\] CPU.registerFile\[24\]\[20\] _07352_ VGND VGND
+ VPWR VPWR _08011_ sky130_fd_sc_hd__mux2_1
X_18115_ net178 _02395_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_16927__7 clknet_1_1__leaf__07220_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__inv_2
XFILLER_0_5_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15327_ _05049_ VGND VGND VPWR VPWR _02826_ sky130_fd_sc_hd__buf_4
XFILLER_0_136_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12539_ net2502 _04779_ _07085_ VGND VGND VPWR VPWR _07092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14438__568 clknet_1_0__leaf__02659_ VGND VGND VPWR VPWR net600 sky130_fd_sc_hd__inv_2
XFILLER_0_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18046_ net1219 _02326_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15258_ _08407_ VGND VGND VPWR VPWR _02757_ sky130_fd_sc_hd__buf_2
XFILLER_0_10_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09750_ mapped_spi_ram.rcv_data\[8\] net16 _04690_ mapped_spi_flash.rcv_data\[8\]
+ VGND VGND VPWR VPWR _05439_ sky130_fd_sc_hd__a22o_2
X_08701_ _04284_ CPU.aluIn1\[4\] VGND VGND VPWR VPWR _04421_ sky130_fd_sc_hd__and2b_1
X_09681_ _04417_ _04806_ _04211_ _04287_ VGND VGND VPWR VPWR _05373_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_107_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14904__988 clknet_1_1__leaf__02705_ VGND VGND VPWR VPWR net1020 sky130_fd_sc_hd__inv_2
X_08632_ CPU.aluIn1\[25\] _04233_ VGND VGND VPWR VPWR _04352_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14603__716 clknet_1_0__leaf__02676_ VGND VGND VPWR VPWR net748 sky130_fd_sc_hd__inv_2
X_08563_ _04282_ VGND VGND VPWR VPWR _04283_ sky130_fd_sc_hd__inv_2
X_15118__1149 clknet_1_0__leaf__02724_ VGND VGND VPWR VPWR net1181 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_120_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08494_ _04213_ VGND VGND VPWR VPWR _04214_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14796__890 clknet_1_0__leaf__02695_ VGND VGND VPWR VPWR net922 sky130_fd_sc_hd__inv_2
XFILLER_0_146_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_804 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09115_ CPU.PC\[20\] _04826_ VGND VGND VPWR VPWR _04827_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09046_ CPU.Bimm\[6\] _04498_ _04760_ VGND VGND VPWR VPWR _04761_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_135_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold440 CPU.registerFile\[2\]\[3\] VGND VGND VPWR VPWR net1681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold451 CPU.registerFile\[28\]\[23\] VGND VGND VPWR VPWR net1692 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 CPU.registerFile\[12\]\[20\] VGND VGND VPWR VPWR net1703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 CPU.registerFile\[14\]\[16\] VGND VGND VPWR VPWR net1714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 CPU.registerFile\[6\]\[15\] VGND VGND VPWR VPWR net1725 sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 CPU.registerFile\[27\]\[2\] VGND VGND VPWR VPWR net1736 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09948_ _05503_ net2329 _05559_ VGND VGND VPWR VPWR _05566_ sky130_fd_sc_hd__mux2_1
X_15069__1134 clknet_1_1__leaf__02723_ VGND VGND VPWR VPWR net1166 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_5_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09879_ _05520_ net2039 _05512_ VGND VGND VPWR VPWR _05521_ sky130_fd_sc_hd__mux2_1
Xhold1140 CPU.registerFile\[10\]\[11\] VGND VGND VPWR VPWR net2381 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1151 CPU.registerFile\[8\]\[13\] VGND VGND VPWR VPWR net2392 sky130_fd_sc_hd__dlygate4sd3_1
X_11910_ net2416 _05689_ _06711_ VGND VGND VPWR VPWR _06721_ sky130_fd_sc_hd__mux2_1
Xhold1162 CPU.registerFile\[14\]\[10\] VGND VGND VPWR VPWR net2403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1173 CPU.registerFile\[18\]\[14\] VGND VGND VPWR VPWR net2414 sky130_fd_sc_hd__dlygate4sd3_1
X_12890_ _07330_ _07331_ VGND VGND VPWR VPWR _07332_ sky130_fd_sc_hd__or2_1
X_14879__965 clknet_1_0__leaf__02703_ VGND VGND VPWR VPWR net997 sky130_fd_sc_hd__inv_2
Xhold1184 mapped_spi_flash.cmd_addr\[22\] VGND VGND VPWR VPWR net2425 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1195 CPU.registerFile\[4\]\[19\] VGND VGND VPWR VPWR net2436 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_302 _07404_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_313 _07914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11841_ _06684_ VGND VGND VPWR VPWR _01647_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_324 _07914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_335 _02887_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_346 _05338_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_357 _07268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_368 _03631_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11772_ _04933_ net2087 _06639_ VGND VGND VPWR VPWR _06648_ sky130_fd_sc_hd__mux2_1
XANTENNA_379 _07530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13511_ _07369_ _07933_ _07935_ _07570_ VGND VGND VPWR VPWR _07936_ sky130_fd_sc_hd__a211o_1
XFILLER_0_83_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10723_ _05530_ net1860 _06045_ VGND VGND VPWR VPWR _06055_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_155_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_138_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16230_ _02797_ _03702_ _03703_ _03704_ _02807_ VGND VGND VPWR VPWR _03705_ sky130_fd_sc_hd__a221o_1
X_13442_ _07653_ _07867_ _07868_ VGND VGND VPWR VPWR _07869_ sky130_fd_sc_hd__o21ai_1
X_10654_ net1337 _06012_ _06013_ VGND VGND VPWR VPWR _02165_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_24_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13373_ CPU.registerFile\[6\]\[14\] CPU.registerFile\[7\]\[14\] _07641_ VGND VGND
+ VPWR VPWR _07802_ sky130_fd_sc_hd__mux2_1
X_16161_ CPU.registerFile\[9\]\[22\] CPU.registerFile\[13\]\[22\] _02887_ VGND VGND
+ VPWR VPWR _03638_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10585_ mapped_spi_flash.rcv_data\[28\] _05970_ VGND VGND VPWR VPWR _05974_ sky130_fd_sc_hd__or2_1
Xclkload18 clknet_leaf_0_clk VGND VGND VPWR VPWR clkload18/Y sky130_fd_sc_hd__inv_8
Xclkload29 clknet_1_0__leaf__03964_ VGND VGND VPWR VPWR clkload29/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_58_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_883 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12324_ _06978_ VGND VGND VPWR VPWR _01423_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16092_ CPU.registerFile\[21\]\[20\] CPU.registerFile\[23\]\[20\] _02769_ VGND VGND
+ VPWR VPWR _03571_ sky130_fd_sc_hd__mux2_1
X_15161__1188 clknet_1_1__leaf__02746_ VGND VGND VPWR VPWR net1220 sky130_fd_sc_hd__inv_2
X_12255_ CPU.aluReg\[16\] CPU.aluReg\[14\] _06906_ VGND VGND VPWR VPWR _06926_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11206_ _05535_ net2415 _06310_ VGND VGND VPWR VPWR _06312_ sky130_fd_sc_hd__mux2_1
X_12186_ CPU.aluReg\[31\] CPU.Bimm\[10\] _06872_ VGND VGND VPWR VPWR _06873_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_71_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11137_ _06275_ VGND VGND VPWR VPWR _01945_ sky130_fd_sc_hd__clkbuf_1
X_16994_ clknet_leaf_28_clk _01320_ VGND VGND VPWR VPWR CPU.rs2\[25\] sky130_fd_sc_hd__dfxtp_1
X_11068_ _06238_ VGND VGND VPWR VPWR _01977_ sky130_fd_sc_hd__clkbuf_1
X_15945_ _05384_ _03425_ _03428_ VGND VGND VPWR VPWR _03429_ sky130_fd_sc_hd__or3_1
XFILLER_0_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10019_ net2354 _04798_ _05596_ VGND VGND VPWR VPWR _05604_ sky130_fd_sc_hd__mux2_1
X_15876_ _02926_ _03360_ _03361_ VGND VGND VPWR VPWR _03362_ sky130_fd_sc_hd__o21a_1
X_17615_ net804 _01903_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17546_ net735 _01834_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13709_ CPU.registerFile\[15\]\[24\] _07236_ _07239_ CPU.registerFile\[11\]\[24\]
+ _07820_ VGND VGND VPWR VPWR _08128_ sky130_fd_sc_hd__o221a_1
X_17477_ net666 _01765_ VGND VGND VPWR VPWR mapped_spi_flash.div_counter\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16428_ CPU.registerFile\[15\]\[30\] CPU.registerFile\[11\]\[30\] _02849_ VGND VGND
+ VPWR VPWR _03897_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_4_Left_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16359_ CPU.registerFile\[14\]\[28\] CPU.registerFile\[10\]\[28\] _02787_ VGND VGND
+ VPWR VPWR _03830_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14371__508 clknet_1_1__leaf__02652_ VGND VGND VPWR VPWR net540 sky130_fd_sc_hd__inv_2
X_18029_ net1202 _02309_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09802_ net2461 _05150_ _05463_ VGND VGND VPWR VPWR _05472_ sky130_fd_sc_hd__mux2_1
X_09733_ CPU.aluReg\[1\] _04219_ _05421_ _05422_ VGND VGND VPWR VPWR _05423_ sky130_fd_sc_hd__a211o_1
X_09664_ _04974_ _05345_ _05347_ _04955_ _05356_ VGND VGND VPWR VPWR _05357_ sky130_fd_sc_hd__o221ai_2
X_08615_ CPU.aluIn1\[16\] _04254_ _04334_ VGND VGND VPWR VPWR _04335_ sky130_fd_sc_hd__a21oi_2
X_09595_ _05288_ _05289_ VGND VGND VPWR VPWR _05290_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08546_ _04264_ _04265_ VGND VGND VPWR VPWR _04266_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08477_ CPU.instr\[3\] CPU.instr\[4\] CPU.instr\[6\] VGND VGND VPWR VPWR _04197_
+ sky130_fd_sc_hd__or3b_4
XFILLER_0_9_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_792 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10370_ _05547_ net1964 _05799_ VGND VGND VPWR VPWR _05807_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_149_Right_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_150_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_522 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09029_ _04504_ _04744_ _04655_ VGND VGND VPWR VPWR _04745_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_131_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12040_ _04780_ net1829 _06783_ VGND VGND VPWR VPWR _06790_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold270 net6 VGND VGND VPWR VPWR net1511 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold281 mapped_spi_flash.rcv_bitcount\[4\] VGND VGND VPWR VPWR net1522 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 CPU.rs2\[15\] VGND VGND VPWR VPWR net1533 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_148_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15730_ CPU.registerFile\[19\]\[9\] CPU.registerFile\[17\]\[9\] _02874_ VGND VGND
+ VPWR VPWR _03220_ sky130_fd_sc_hd__mux2_1
X_12942_ _07283_ VGND VGND VPWR VPWR _07383_ sky130_fd_sc_hd__clkbuf_8
X_14467__594 clknet_1_0__leaf__02662_ VGND VGND VPWR VPWR net626 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_29_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15661_ CPU.registerFile\[22\]\[7\] CPU.registerFile\[23\]\[7\] _02828_ VGND VGND
+ VPWR VPWR _03153_ sky130_fd_sc_hd__mux2_1
XANTENNA_110 _05406_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12873_ _07314_ VGND VGND VPWR VPWR _07315_ sky130_fd_sc_hd__buf_8
XANTENNA_121 _05526_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_132 _05551_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17400_ net589 _01688_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_bitcount\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_143 _07231_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11824_ net2249 _05668_ _06675_ VGND VGND VPWR VPWR _06676_ sky130_fd_sc_hd__mux2_1
XANTENNA_154 _07271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15592_ CPU.registerFile\[8\]\[6\] _02763_ _02764_ _03084_ VGND VGND VPWR VPWR _03085_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_165 _07325_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_176 _07476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17331_ net520 _01619_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_187 _07841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_198 _07841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11755_ _06638_ VGND VGND VPWR VPWR _06639_ sky130_fd_sc_hd__buf_4
XFILLER_0_154_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10706_ _06046_ VGND VGND VPWR VPWR _02147_ sky130_fd_sc_hd__clkbuf_1
X_17262_ net452 _01550_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11686_ mapped_spi_ram.rcv_data\[17\] _06588_ VGND VGND VPWR VPWR _06596_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16213_ CPU.registerFile\[25\]\[23\] CPU.registerFile\[29\]\[23\] _02798_ VGND VGND
+ VPWR VPWR _03689_ sky130_fd_sc_hd__mux2_1
X_13425_ CPU.registerFile\[13\]\[15\] _07361_ _07521_ CPU.registerFile\[9\]\[15\]
+ _07285_ VGND VGND VPWR VPWR _07853_ sky130_fd_sc_hd__o221a_1
X_17193_ clknet_leaf_25_clk _01481_ VGND VGND VPWR VPWR CPU.Iimm\[3\] sky130_fd_sc_hd__dfxtp_2
X_10637_ net1395 _05994_ VGND VGND VPWR VPWR _06003_ sky130_fd_sc_hd__or2_1
Xclkload107 clknet_1_1__leaf__08358_ VGND VGND VPWR VPWR clkload107/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload118 clknet_1_0__leaf__07220_ VGND VGND VPWR VPWR clkload118/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_3_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16144_ _03618_ _03619_ _03621_ _02812_ VGND VGND VPWR VPWR _03622_ sky130_fd_sc_hd__o22a_2
X_13356_ CPU.registerFile\[18\]\[13\] CPU.registerFile\[22\]\[13\] _07785_ VGND VGND
+ VPWR VPWR _07786_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_116_Right_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10568_ _05952_ _05950_ mapped_spi_flash.snd_bitcount\[0\] VGND VGND VPWR VPWR _05961_
+ sky130_fd_sc_hd__mux2_1
X_14632__742 clknet_1_1__leaf__02679_ VGND VGND VPWR VPWR net774 sky130_fd_sc_hd__inv_2
XFILLER_0_122_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12307_ net2435 _06965_ _06861_ VGND VGND VPWR VPWR _06966_ sky130_fd_sc_hd__mux2_1
X_16075_ CPU.registerFile\[25\]\[19\] CPU.registerFile\[29\]\[19\] _03254_ VGND VGND
+ VPWR VPWR _03555_ sky130_fd_sc_hd__mux2_1
X_15117__1148 clknet_1_0__leaf__02724_ VGND VGND VPWR VPWR net1180 sky130_fd_sc_hd__inv_2
X_13287_ CPU.registerFile\[1\]\[11\] _07387_ _07718_ _07231_ VGND VGND VPWR VPWR _07719_
+ sky130_fd_sc_hd__a211o_1
X_10499_ _05886_ _05906_ VGND VGND VPWR VPWR _05907_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12238_ CPU.aluReg\[20\] CPU.aluReg\[18\] _06906_ VGND VGND VPWR VPWR _06913_ sky130_fd_sc_hd__mux2_1
X_12169_ _04589_ _06860_ VGND VGND VPWR VPWR _06861_ sky130_fd_sc_hd__nor2_4
X_16977_ clknet_leaf_26_clk _01303_ VGND VGND VPWR VPWR CPU.rs2\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_88_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15928_ _08401_ _03408_ _03411_ _02844_ VGND VGND VPWR VPWR _03412_ sky130_fd_sc_hd__o211a_1
X_15859_ _02911_ _03342_ _03344_ _02794_ VGND VGND VPWR VPWR _03345_ sky130_fd_sc_hd__a211o_1
X_09380_ _04899_ _05084_ VGND VGND VPWR VPWR _05085_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17529_ net718 _01817_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[11\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_49_Left_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14715__817 clknet_1_1__leaf__02687_ VGND VGND VPWR VPWR net849 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_15_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15068__1133 clknet_1_1__leaf__02723_ VGND VGND VPWR VPWR net1165 sky130_fd_sc_hd__inv_2
XFILLER_0_117_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14295__439 clknet_1_1__leaf__08462_ VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__inv_2
XFILLER_0_144_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_58_Left_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14761__859 clknet_1_1__leaf__02691_ VGND VGND VPWR VPWR net891 sky130_fd_sc_hd__inv_2
X_09716_ _05405_ VGND VGND VPWR VPWR _05406_ sky130_fd_sc_hd__buf_4
XFILLER_0_69_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16521__189 clknet_1_1__leaf__03963_ VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__inv_2
X_09647_ mapped_spi_flash.rcv_data\[28\] _04784_ _05339_ VGND VGND VPWR VPWR _05340_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_143_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15160__1187 clknet_1_1__leaf__02746_ VGND VGND VPWR VPWR net1219 sky130_fd_sc_hd__inv_2
X_09578_ net1894 _05273_ _05189_ VGND VGND VPWR VPWR _05274_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_67_Left_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08529_ CPU.rs2\[18\] _04200_ _04205_ VGND VGND VPWR VPWR _04249_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11540_ _06494_ VGND VGND VPWR VPWR _06495_ sky130_fd_sc_hd__buf_2
XFILLER_0_148_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11471_ _06452_ VGND VGND VPWR VPWR _01788_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13210_ CPU.registerFile\[3\]\[9\] _07373_ _07376_ VGND VGND VPWR VPWR _07644_ sky130_fd_sc_hd__o21a_1
X_10422_ net1369 _05841_ _05842_ net1347 _05844_ VGND VGND VPWR VPWR _02228_ sky130_fd_sc_hd__o221a_1
XFILLER_0_150_447 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13141_ _04986_ VGND VGND VPWR VPWR _07577_ sky130_fd_sc_hd__buf_4
XFILLER_0_131_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10353_ _05530_ net2150 _05788_ VGND VGND VPWR VPWR _05798_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_76_Left_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13072_ _07508_ _07509_ _07315_ VGND VGND VPWR VPWR _07510_ sky130_fd_sc_hd__mux2_1
X_10284_ _05530_ net2014 _05751_ VGND VGND VPWR VPWR _05761_ sky130_fd_sc_hd__mux2_1
X_12023_ _06780_ VGND VGND VPWR VPWR _01561_ sky130_fd_sc_hd__clkbuf_1
X_16900_ _04644_ _06468_ VGND VGND VPWR VPWR _04177_ sky130_fd_sc_hd__and2_1
X_17880_ net1069 _02164_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_bitcount\[5\] sky130_fd_sc_hd__dfxtp_1
X_16831_ per_uart.uart0.tx_bitcount\[2\] per_uart.uart0.tx_bitcount\[1\] per_uart.uart0.tx_bitcount\[0\]
+ VGND VGND VPWR VPWR _04131_ sky130_fd_sc_hd__and3_1
X_16762_ _08379_ _04926_ _05062_ _08454_ VGND VGND VPWR VPWR _04078_ sky130_fd_sc_hd__or4b_1
X_15713_ CPU.registerFile\[6\]\[9\] CPU.registerFile\[7\]\[9\] _02870_ VGND VGND VPWR
+ VPWR _03203_ sky130_fd_sc_hd__mux2_1
X_12925_ _07364_ _07365_ VGND VGND VPWR VPWR _07366_ sky130_fd_sc_hd__or2_1
X_16693_ _04001_ _04017_ _04018_ _04019_ _07123_ VGND VGND VPWR VPWR _04020_ sky130_fd_sc_hd__o311a_1
X_16496__166 clknet_1_0__leaf__02756_ VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_66_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_85_Left_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15644_ CPU.registerFile\[25\]\[7\] _02802_ _02803_ VGND VGND VPWR VPWR _03136_ sky130_fd_sc_hd__o21a_1
X_12856_ _07296_ _07298_ VGND VGND VPWR VPWR _07299_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11807_ _06666_ VGND VGND VPWR VPWR _01663_ sky130_fd_sc_hd__clkbuf_1
X_18363_ clknet_leaf_9_clk _02641_ VGND VGND VPWR VPWR per_uart.d_in_uart\[3\] sky130_fd_sc_hd__dfxtp_1
X_15575_ _02834_ VGND VGND VPWR VPWR _03069_ sky130_fd_sc_hd__clkbuf_4
X_12787_ _04814_ VGND VGND VPWR VPWR _07230_ sky130_fd_sc_hd__clkbuf_4
X_17314_ net503 _01602_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18294_ net127 _02574_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_11738_ _06624_ net1755 _06627_ VGND VGND VPWR VPWR _06628_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_731 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17245_ net435 _01533_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11669_ net1434 _06577_ VGND VGND VPWR VPWR _06586_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13408_ _07260_ _07835_ VGND VGND VPWR VPWR _07836_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17176_ clknet_leaf_12_clk _01464_ VGND VGND VPWR VPWR CPU.instr\[6\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_94_Left_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16127_ CPU.registerFile\[9\]\[21\] _02802_ _03125_ VGND VGND VPWR VPWR _03605_ sky130_fd_sc_hd__o21a_1
X_13339_ CPU.registerFile\[14\]\[13\] CPU.registerFile\[10\]\[13\] _04936_ VGND VGND
+ VPWR VPWR _07769_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16058_ CPU.registerFile\[22\]\[19\] _08399_ VGND VGND VPWR VPWR _03538_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__02696_ clknet_0__02696_ VGND VGND VPWR VPWR clknet_1_1__leaf__02696_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_94_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__07223_ clknet_0__07223_ VGND VGND VPWR VPWR clknet_1_1__leaf__07223_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_110_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_889 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08880_ _04558_ _04561_ _04590_ VGND VGND VPWR VPWR _04600_ sky130_fd_sc_hd__o21a_1
XFILLER_0_138_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14483__609 clknet_1_0__leaf__02663_ VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__inv_2
X_09501_ _04266_ _04402_ _04429_ VGND VGND VPWR VPWR _05200_ sky130_fd_sc_hd__nor3_1
XFILLER_0_154_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09432_ _04216_ _04208_ VGND VGND VPWR VPWR _05134_ sky130_fd_sc_hd__nand2_2
XFILLER_0_154_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09363_ _04594_ _04599_ _04613_ VGND VGND VPWR VPWR _05068_ sky130_fd_sc_hd__nor3_1
XFILLER_0_157_580 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14303__446 clknet_1_1__leaf__08463_ VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__inv_2
X_09294_ _05001_ _05002_ VGND VGND VPWR VPWR _05003_ sky130_fd_sc_hd__or2_1
XANTENNA_10 _02842_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_21 _02940_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_32 _03077_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 _04483_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_54 _04971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_65 _05090_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 _05169_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_87 _05284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_98 _05359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_924 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_132_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_145_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__08430_ clknet_0__08430_ VGND VGND VPWR VPWR clknet_1_0__leaf__08430_
+ sky130_fd_sc_hd__clkbuf_16
X_10971_ net1632 _05685_ _06179_ VGND VGND VPWR VPWR _06187_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__08361_ clknet_0__08361_ VGND VGND VPWR VPWR clknet_1_0__leaf__08361_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_39_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12710_ net1465 _07191_ VGND VGND VPWR VPWR _07192_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_39_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13690_ _08105_ _08106_ _08107_ _08109_ _04814_ VGND VGND VPWR VPWR _08110_ sky130_fd_sc_hd__a221o_1
X_15116__1147 clknet_1_0__leaf__02724_ VGND VGND VPWR VPWR net1179 sky130_fd_sc_hd__inv_2
XFILLER_0_66_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12641_ CPU.cycles\[9\] _07144_ VGND VGND VPWR VPWR _07146_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14579__695 clknet_1_1__leaf__02673_ VGND VGND VPWR VPWR net727 sky130_fd_sc_hd__inv_2
X_15360_ _02758_ VGND VGND VPWR VPWR _02858_ sky130_fd_sc_hd__clkbuf_8
X_12572_ _07109_ VGND VGND VPWR VPWR _01273_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11523_ net1334 mapped_spi_ram.snd_bitcount\[2\] _06483_ _06484_ VGND VGND VPWR VPWR
+ _06485_ sky130_fd_sc_hd__nor4_1
X_15291_ _05070_ VGND VGND VPWR VPWR _02790_ sky130_fd_sc_hd__buf_4
XFILLER_0_135_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17030_ net288 _01352_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_11454_ _06443_ VGND VGND VPWR VPWR _01796_ sky130_fd_sc_hd__clkbuf_1
X_10405_ mapped_spi_flash.cmd_addr\[28\] _05825_ _05827_ mapped_spi_flash.cmd_addr\[29\]
+ VGND VGND VPWR VPWR _05833_ sky130_fd_sc_hd__a22o_1
X_11385_ _05509_ net2221 _06397_ VGND VGND VPWR VPWR _06407_ sky130_fd_sc_hd__mux2_1
X_14173_ CPU.Bimm\[9\] _04710_ _08413_ VGND VGND VPWR VPWR _08424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13124_ CPU.registerFile\[31\]\[6\] _07347_ _07348_ CPU.registerFile\[27\]\[6\] _07345_
+ VGND VGND VPWR VPWR _07561_ sky130_fd_sc_hd__o221a_1
X_10336_ _05789_ VGND VGND VPWR VPWR _02260_ sky130_fd_sc_hd__clkbuf_1
X_13055_ CPU.registerFile\[15\]\[4\] _07402_ _07420_ CPU.registerFile\[11\]\[4\] _07483_
+ VGND VGND VPWR VPWR _07494_ sky130_fd_sc_hd__o221a_1
X_10267_ _05752_ VGND VGND VPWR VPWR _02307_ sky130_fd_sc_hd__clkbuf_1
X_17932_ net1121 _02216_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[12\] sky130_fd_sc_hd__dfxtp_1
X_12006_ _05230_ net2357 _06769_ VGND VGND VPWR VPWR _06772_ sky130_fd_sc_hd__mux2_1
X_17863_ net1052 _02147_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_10198_ _05149_ VGND VGND VPWR VPWR _05708_ sky130_fd_sc_hd__clkbuf_4
X_14744__843 clknet_1_0__leaf__02690_ VGND VGND VPWR VPWR net875 sky130_fd_sc_hd__inv_2
X_15067__1132 clknet_1_0__leaf__02723_ VGND VGND VPWR VPWR net1164 sky130_fd_sc_hd__inv_2
X_16814_ _08355_ _07196_ _04117_ _04118_ per_uart.uart0.tx_count16\[1\] VGND VGND
+ VPWR VPWR _04119_ sky130_fd_sc_hd__a32o_1
X_17794_ net983 _02078_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_16504__173 clknet_1_1__leaf__03962_ VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__inv_2
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16745_ _03995_ _05118_ _07132_ VGND VGND VPWR VPWR _04064_ sky130_fd_sc_hd__o21ai_1
X_12908_ CPU.registerFile\[29\]\[1\] _07347_ _07348_ CPU.registerFile\[25\]\[1\] _07349_
+ VGND VGND VPWR VPWR _07350_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_17_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16676_ _08436_ _08459_ _05345_ VGND VGND VPWR VPWR _04005_ sky130_fd_sc_hd__a21o_1
X_13888_ _07330_ _08300_ VGND VGND VPWR VPWR _08301_ sky130_fd_sc_hd__or2_1
XFILLER_0_158_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15627_ CPU.registerFile\[12\]\[7\] _03118_ VGND VGND VPWR VPWR _03119_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12839_ _07281_ VGND VGND VPWR VPWR _07282_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_158_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18346_ clknet_leaf_1_clk _02626_ VGND VGND VPWR VPWR per_uart.uart0.rx_count16\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_15558_ CPU.registerFile\[29\]\[5\] _02800_ VGND VGND VPWR VPWR _03052_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18277_ net110 _02557_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_14790__885 clknet_1_1__leaf__02694_ VGND VGND VPWR VPWR net917 sky130_fd_sc_hd__inv_2
X_15489_ _05361_ _02984_ VGND VGND VPWR VPWR _02985_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17228_ net418 _01516_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[21\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03966_ _03966_ VGND VGND VPWR VPWR clknet_0__03966_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold803 CPU.registerFile\[4\]\[18\] VGND VGND VPWR VPWR net2044 sky130_fd_sc_hd__dlygate4sd3_1
X_17159_ net383 _01447_ VGND VGND VPWR VPWR CPU.aluReg\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_678 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold814 CPU.registerFile\[24\]\[18\] VGND VGND VPWR VPWR net2055 sky130_fd_sc_hd__dlygate4sd3_1
Xhold825 CPU.registerFile\[12\]\[22\] VGND VGND VPWR VPWR net2066 sky130_fd_sc_hd__dlygate4sd3_1
Xhold836 CPU.registerFile\[12\]\[16\] VGND VGND VPWR VPWR net2077 sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 CPU.registerFile\[14\]\[7\] VGND VGND VPWR VPWR net2088 sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 CPU.registerFile\[22\]\[2\] VGND VGND VPWR VPWR net2099 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__02748_ clknet_0__02748_ VGND VGND VPWR VPWR clknet_1_1__leaf__02748_
+ sky130_fd_sc_hd__clkbuf_16
X_09981_ _05583_ VGND VGND VPWR VPWR _02456_ sky130_fd_sc_hd__clkbuf_1
Xhold869 CPU.registerFile\[28\]\[21\] VGND VGND VPWR VPWR net2110 sky130_fd_sc_hd__dlygate4sd3_1
X_14827__918 clknet_1_0__leaf__02698_ VGND VGND VPWR VPWR net950 sky130_fd_sc_hd__inv_2
X_08932_ _04484_ _04622_ _04651_ _04483_ VGND VGND VPWR VPWR _04652_ sky130_fd_sc_hd__a211o_1
Xclkbuf_1_1__f__02679_ clknet_0__02679_ VGND VGND VPWR VPWR clknet_1_1__leaf__02679_
+ sky130_fd_sc_hd__clkbuf_16
X_08863_ CPU.aluIn1\[21\] _04495_ VGND VGND VPWR VPWR _04583_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08794_ CPU.aluIn1\[8\] CPU.Bimm\[8\] VGND VGND VPWR VPWR _04514_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09415_ _04437_ _04328_ VGND VGND VPWR VPWR _05118_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_832 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09346_ CPU.Jimm\[17\] _04812_ _04989_ CPU.cycles\[17\] VGND VGND VPWR VPWR _05052_
+ sky130_fd_sc_hd__a22o_1
X_15210__121 clknet_1_1__leaf__02752_ VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__inv_2
XFILLER_0_75_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09277_ net14 VGND VGND VPWR VPWR _04986_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_133_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11170_ _05499_ net2295 _06288_ VGND VGND VPWR VPWR _06293_ sky130_fd_sc_hd__mux2_1
X_10121_ _05658_ VGND VGND VPWR VPWR _02359_ sky130_fd_sc_hd__clkbuf_1
X_10052_ _05621_ VGND VGND VPWR VPWR _02391_ sky130_fd_sc_hd__clkbuf_1
X_13811_ _07291_ _08226_ VGND VGND VPWR VPWR _08227_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_3_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13742_ CPU.registerFile\[23\]\[25\] _07414_ _08159_ _07621_ _04648_ VGND VGND VPWR
+ VPWR _08160_ sky130_fd_sc_hd__o221a_1
X_10954_ _06177_ VGND VGND VPWR VPWR _02030_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16461_ CPU.registerFile\[1\]\[31\] _03228_ _03928_ _02818_ VGND VGND VPWR VPWR _03929_
+ sky130_fd_sc_hd__a22o_1
X_13673_ CPU.registerFile\[23\]\[23\] _07382_ _08092_ _07818_ VGND VGND VPWR VPWR
+ _08093_ sky130_fd_sc_hd__o22a_1
X_10885_ _06140_ VGND VGND VPWR VPWR _02062_ sky130_fd_sc_hd__clkbuf_1
X_18200_ net231 _02480_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[2\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__02699_ clknet_0__02699_ VGND VGND VPWR VPWR clknet_1_0__leaf__02699_
+ sky130_fd_sc_hd__clkbuf_16
X_15412_ _02907_ _02908_ _02875_ VGND VGND VPWR VPWR _02909_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_158_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12624_ CPU.cycles\[0\] CPU.cycles\[1\] CPU.cycles\[2\] VGND VGND VPWR VPWR _07136_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_109_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_158_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16392_ CPU.aluIn1\[28\] _07358_ _03862_ _03632_ VGND VGND VPWR VPWR _02442_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_158_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__07226_ clknet_0__07226_ VGND VGND VPWR VPWR clknet_1_0__leaf__07226_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_26_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18131_ net194 _02411_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15343_ _02838_ _02841_ _02809_ VGND VGND VPWR VPWR _02842_ sky130_fd_sc_hd__a21oi_4
X_12555_ _07100_ VGND VGND VPWR VPWR _01281_ sky130_fd_sc_hd__clkbuf_1
X_18062_ net1235 _02342_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_11506_ _06471_ _06472_ VGND VGND VPWR VPWR _06473_ sky130_fd_sc_hd__or2_1
X_15274_ _02772_ VGND VGND VPWR VPWR _02773_ sky130_fd_sc_hd__clkbuf_8
X_12486_ net1745 _05698_ _07060_ VGND VGND VPWR VPWR _07064_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17013_ net271 _01335_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11437_ _05493_ net2255 _06433_ VGND VGND VPWR VPWR _06435_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__02702_ _02702_ VGND VGND VPWR VPWR clknet_0__02702_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14156_ CPU.Iimm\[1\] _07380_ _08413_ VGND VGND VPWR VPWR _08415_ sky130_fd_sc_hd__mux2_1
X_11368_ _06398_ VGND VGND VPWR VPWR _01837_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ CPU.registerFile\[7\]\[6\] _07262_ _07543_ _07265_ VGND VGND VPWR VPWR _07544_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_91_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10319_ _05780_ VGND VGND VPWR VPWR _02268_ sky130_fd_sc_hd__clkbuf_1
X_14087_ _04291_ _07134_ VGND VGND VPWR VPWR _08369_ sky130_fd_sc_hd__nor2_1
X_11299_ _06361_ VGND VGND VPWR VPWR _01869_ sky130_fd_sc_hd__clkbuf_1
X_14332__472 clknet_1_0__leaf__08466_ VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__inv_2
X_13038_ CPU.registerFile\[28\]\[4\] CPU.registerFile\[24\]\[4\] _07476_ VGND VGND
+ VPWR VPWR _07477_ sky130_fd_sc_hd__mux2_1
X_17915_ net1104 _02199_ VGND VGND VPWR VPWR mapped_spi_flash.snd_bitcount\[1\] sky130_fd_sc_hd__dfxtp_1
X_13970__254 clknet_1_1__leaf__08357_ VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__inv_2
X_17846_ net1035 _02130_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_17777_ net966 _02061_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_754 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16728_ _03991_ net1623 VGND VGND VPWR VPWR _04049_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16659_ _08455_ VGND VGND VPWR VPWR _03990_ sky130_fd_sc_hd__buf_2
X_09200_ CPU.PC\[23\] _04911_ VGND VGND VPWR VPWR _04912_ sky130_fd_sc_hd__xor2_1
XFILLER_0_56_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09131_ CPU.PC\[16\] _04842_ VGND VGND VPWR VPWR _04843_ sky130_fd_sc_hd__and2_1
X_18329_ clknet_leaf_6_clk _02609_ VGND VGND VPWR VPWR per_uart.uart0.tx_count16\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09062_ mapped_spi_ram.rcv_data\[1\] _04689_ _04691_ mapped_spi_flash.rcv_data\[1\]
+ VGND VGND VPWR VPWR _04776_ sky130_fd_sc_hd__a22o_2
XFILLER_0_72_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12773__222 clknet_1_0__leaf__07225_ VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__inv_2
XFILLER_0_25_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold600 CPU.registerFile\[27\]\[4\] VGND VGND VPWR VPWR net1841 sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 CPU.registerFile\[30\]\[16\] VGND VGND VPWR VPWR net1852 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold622 CPU.registerFile\[29\]\[16\] VGND VGND VPWR VPWR net1863 sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 CPU.registerFile\[3\]\[27\] VGND VGND VPWR VPWR net1874 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14415__547 clknet_1_0__leaf__02657_ VGND VGND VPWR VPWR net579 sky130_fd_sc_hd__inv_2
Xhold644 CPU.registerFile\[22\]\[13\] VGND VGND VPWR VPWR net1885 sky130_fd_sc_hd__dlygate4sd3_1
Xhold655 CPU.registerFile\[30\]\[14\] VGND VGND VPWR VPWR net1896 sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 CPU.registerFile\[17\]\[28\] VGND VGND VPWR VPWR net1907 sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 CPU.registerFile\[30\]\[31\] VGND VGND VPWR VPWR net1918 sky130_fd_sc_hd__dlygate4sd3_1
X_15115__1146 clknet_1_1__leaf__02724_ VGND VGND VPWR VPWR net1178 sky130_fd_sc_hd__inv_2
Xhold688 CPU.registerFile\[3\]\[2\] VGND VGND VPWR VPWR net1929 sky130_fd_sc_hd__dlygate4sd3_1
X_09964_ _05574_ VGND VGND VPWR VPWR _02464_ sky130_fd_sc_hd__clkbuf_1
Xhold699 CPU.registerFile\[23\]\[26\] VGND VGND VPWR VPWR net1940 sky130_fd_sc_hd__dlygate4sd3_1
X_08915_ CPU.PC\[4\] _04598_ _04633_ _04634_ VGND VGND VPWR VPWR _04635_ sky130_fd_sc_hd__a22oi_4
X_09895_ _05531_ VGND VGND VPWR VPWR _02490_ sky130_fd_sc_hd__clkbuf_1
Xhold1300 net12 VGND VGND VPWR VPWR net2541 sky130_fd_sc_hd__dlygate4sd3_1
X_08846_ CPU.aluIn1\[18\] _04494_ VGND VGND VPWR VPWR _04566_ sky130_fd_sc_hd__nand2_1
X_08777_ net1274 CPU.instr\[2\] _04293_ VGND VGND VPWR VPWR _04497_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_0_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14461__589 clknet_1_1__leaf__02661_ VGND VGND VPWR VPWR net621 sky130_fd_sc_hd__inv_2
XFILLER_0_95_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_40_Left_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_662 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10670_ net1346 _06018_ _06022_ _06025_ VGND VGND VPWR VPWR _02162_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09329_ _04388_ _04443_ VGND VGND VPWR VPWR _05036_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclone33 net1275 VGND VGND VPWR VPWR net1274 sky130_fd_sc_hd__clkbuf_16
X_12340_ _06986_ VGND VGND VPWR VPWR _01415_ sky130_fd_sc_hd__clkbuf_1
X_15066__1131 clknet_1_0__leaf__02723_ VGND VGND VPWR VPWR net1163 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_153_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12271_ _06938_ VGND VGND VPWR VPWR _01436_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11222_ _05551_ net2099 _06310_ VGND VGND VPWR VPWR _06320_ sky130_fd_sc_hd__mux2_1
X_11153_ _06283_ VGND VGND VPWR VPWR _01937_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_56_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10104_ _05649_ VGND VGND VPWR VPWR _02367_ sky130_fd_sc_hd__clkbuf_1
X_11084_ _06246_ VGND VGND VPWR VPWR _01969_ sky130_fd_sc_hd__clkbuf_1
X_15961_ CPU.registerFile\[27\]\[16\] CPU.registerFile\[31\]\[16\] _03050_ VGND VGND
+ VPWR VPWR _03444_ sky130_fd_sc_hd__mux2_1
X_17700_ net889 _01988_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_10035_ _05612_ VGND VGND VPWR VPWR _02399_ sky130_fd_sc_hd__clkbuf_1
X_15892_ CPU.registerFile\[24\]\[14\] _03130_ _02790_ _03376_ VGND VGND VPWR VPWR
+ _03377_ sky130_fd_sc_hd__o211a_1
X_17631_ net820 _01919_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_17562_ net751 _01850_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_11986_ _06761_ VGND VGND VPWR VPWR _01579_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13725_ CPU.registerFile\[16\]\[25\] CPU.registerFile\[20\]\[25\] _05283_ VGND VGND
+ VPWR VPWR _08143_ sky130_fd_sc_hd__mux2_1
X_10937_ net1585 _05719_ _06165_ VGND VGND VPWR VPWR _06169_ sky130_fd_sc_hd__mux2_1
X_14856__944 clknet_1_1__leaf__02701_ VGND VGND VPWR VPWR net976 sky130_fd_sc_hd__inv_2
XFILLER_0_86_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17493_ net682 _01781_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16444_ CPU.registerFile\[30\]\[30\] CPU.registerFile\[26\]\[30\] _02773_ VGND VGND
+ VPWR VPWR _03913_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13656_ _08072_ _08073_ _08076_ _07250_ _07359_ VGND VGND VPWR VPWR _08077_ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10868_ net2478 _05719_ _06128_ VGND VGND VPWR VPWR _06132_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12607_ CPU.state\[2\] _07120_ VGND VGND VPWR VPWR _07126_ sky130_fd_sc_hd__nand2_1
X_16375_ _02885_ _03843_ _03844_ _03845_ _03022_ VGND VGND VPWR VPWR _03846_ sky130_fd_sc_hd__a221o_1
X_13587_ CPU.registerFile\[29\]\[20\] _07347_ _07348_ CPU.registerFile\[25\]\[20\]
+ _07300_ VGND VGND VPWR VPWR _08010_ sky130_fd_sc_hd__o221a_1
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10799_ _06095_ VGND VGND VPWR VPWR _02103_ sky130_fd_sc_hd__clkbuf_1
X_18114_ net177 _02394_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_15326_ _02812_ _02817_ _02824_ _02809_ VGND VGND VPWR VPWR _02825_ sky130_fd_sc_hd__o211a_1
X_12538_ _07091_ VGND VGND VPWR VPWR _01289_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18045_ net1218 _02325_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_12469_ net1987 _05681_ _07049_ VGND VGND VPWR VPWR _07055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14139_ _08402_ VGND VGND VPWR VPWR _01474_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_120_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08700_ _04407_ _04418_ _04419_ VGND VGND VPWR VPWR _04420_ sky130_fd_sc_hd__o21a_1
X_09680_ CPU.aluIn1\[3\] _04286_ _04214_ _04219_ CPU.aluReg\[3\] VGND VGND VPWR VPWR
+ _05372_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_107_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08631_ _04347_ _04238_ _04348_ _04350_ VGND VGND VPWR VPWR _04351_ sky130_fd_sc_hd__o211a_1
X_17829_ net1018 _02113_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_08562_ _04280_ _04281_ VGND VGND VPWR VPWR _04282_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08493_ CPU.Jimm\[13\] CPU.Jimm\[14\] _04208_ VGND VGND VPWR VPWR _04213_ sky130_fd_sc_hd__and3_1
XFILLER_0_147_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09114_ CPU.Iimm\[0\] _04496_ _04820_ VGND VGND VPWR VPWR _04826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09045_ CPU.cycles\[26\] _04503_ _04757_ _04708_ _04759_ VGND VGND VPWR VPWR _04760_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_135_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold430 CPU.registerFile\[18\]\[25\] VGND VGND VPWR VPWR net1671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 CPU.registerFile\[12\]\[18\] VGND VGND VPWR VPWR net1682 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold452 CPU.registerFile\[30\]\[26\] VGND VGND VPWR VPWR net1693 sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 mapped_spi_flash.rcv_data\[23\] VGND VGND VPWR VPWR net1704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold474 CPU.registerFile\[5\]\[23\] VGND VGND VPWR VPWR net1715 sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 CPU.registerFile\[12\]\[11\] VGND VGND VPWR VPWR net1726 sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 CPU.registerFile\[16\]\[10\] VGND VGND VPWR VPWR net1737 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09947_ _05565_ VGND VGND VPWR VPWR _02472_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_5_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ _05065_ VGND VGND VPWR VPWR _05520_ sky130_fd_sc_hd__buf_6
Xhold1130 CPU.registerFile\[25\]\[3\] VGND VGND VPWR VPWR net2371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1141 CPU.registerFile\[1\]\[14\] VGND VGND VPWR VPWR net2382 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1152 CPU.registerFile\[2\]\[18\] VGND VGND VPWR VPWR net2393 sky130_fd_sc_hd__dlygate4sd3_1
X_08829_ CPU.aluIn1\[11\] CPU.Bimm\[12\] VGND VGND VPWR VPWR _04549_ sky130_fd_sc_hd__or2_1
Xhold1163 CPU.registerFile\[1\]\[2\] VGND VGND VPWR VPWR net2404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1174 CPU.registerFile\[22\]\[10\] VGND VGND VPWR VPWR net2415 sky130_fd_sc_hd__dlygate4sd3_1
X_14014__294 clknet_1_0__leaf__08361_ VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__inv_2
Xhold1185 CPU.registerFile\[23\]\[17\] VGND VGND VPWR VPWR net2426 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1196 CPU.registerFile\[11\]\[29\] VGND VGND VPWR VPWR net2437 sky130_fd_sc_hd__dlygate4sd3_1
X_11840_ CPU.registerFile\[10\]\[23\] _05687_ _06675_ VGND VGND VPWR VPWR _06684_
+ sky130_fd_sc_hd__mux2_1
XANTENNA_303 _07404_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_314 _07914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_325 _07914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_336 _02887_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_347 _05338_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_358 _07268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11771_ _06647_ VGND VGND VPWR VPWR _01680_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_369 _05188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_13510_ CPU.registerFile\[3\]\[18\] _07373_ _07934_ _07376_ VGND VGND VPWR VPWR _07935_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_24_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ _06054_ VGND VGND VPWR VPWR _02139_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_155_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13441_ CPU.registerFile\[21\]\[16\] _07403_ _07404_ CPU.registerFile\[17\]\[16\]
+ _07250_ VGND VGND VPWR VPWR _07868_ sky130_fd_sc_hd__o221a_1
X_10653_ net7 _06012_ _04193_ VGND VGND VPWR VPWR _06013_ sky130_fd_sc_hd__o21a_1
XFILLER_0_24_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16160_ CPU.registerFile\[11\]\[22\] _02895_ _02924_ _03636_ VGND VGND VPWR VPWR
+ _03637_ sky130_fd_sc_hd__o211a_1
X_13372_ _07638_ VGND VGND VPWR VPWR _07801_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10584_ net1483 _05968_ _05973_ _05936_ VGND VGND VPWR VPWR _02195_ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload19 clknet_leaf_2_clk VGND VGND VPWR VPWR clkload19/Y sky130_fd_sc_hd__inv_6
X_15111_ _02742_ VGND VGND VPWR VPWR _02285_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12323_ _04659_ net2160 _06977_ VGND VGND VPWR VPWR _06978_ sky130_fd_sc_hd__mux2_1
X_16091_ _03566_ _03569_ _02858_ VGND VGND VPWR VPWR _03570_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_895 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15042_ clknet_1_1__leaf__02720_ VGND VGND VPWR VPWR _02721_ sky130_fd_sc_hd__buf_1
X_12254_ _06925_ VGND VGND VPWR VPWR _01440_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11205_ _06311_ VGND VGND VPWR VPWR _01913_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_71_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12185_ _04483_ _05134_ VGND VGND VPWR VPWR _06872_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_71_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11136_ net2358 _05712_ _06274_ VGND VGND VPWR VPWR _06275_ sky130_fd_sc_hd__mux2_1
X_16993_ clknet_leaf_21_clk _01319_ VGND VGND VPWR VPWR CPU.rs2\[24\] sky130_fd_sc_hd__dfxtp_1
X_11067_ net1833 _05712_ _06237_ VGND VGND VPWR VPWR _06238_ sky130_fd_sc_hd__mux2_1
X_15944_ _03030_ _03426_ _03427_ _02901_ VGND VGND VPWR VPWR _03428_ sky130_fd_sc_hd__a22o_1
X_10018_ _05603_ VGND VGND VPWR VPWR _02407_ sky130_fd_sc_hd__clkbuf_1
X_15875_ CPU.registerFile\[18\]\[13\] _02832_ _02835_ CPU.registerFile\[19\]\[13\]
+ _03074_ VGND VGND VPWR VPWR _03361_ sky130_fd_sc_hd__o221a_1
X_17614_ net803 _01902_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14444__573 clknet_1_1__leaf__02660_ VGND VGND VPWR VPWR net605 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_102_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17545_ net734 _01833_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11969_ _06752_ VGND VGND VPWR VPWR _01587_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13708_ CPU.registerFile\[14\]\[24\] CPU.registerFile\[10\]\[24\] _07480_ VGND VGND
+ VPWR VPWR _08127_ sky130_fd_sc_hd__mux2_1
X_14182__361 clknet_1_1__leaf__08428_ VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__inv_2
X_15114__1145 clknet_1_1__leaf__02724_ VGND VGND VPWR VPWR net1177 sky130_fd_sc_hd__inv_2
XFILLER_0_46_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17476_ net665 _01764_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16427_ net2497 _07228_ _03877_ _03896_ _06482_ VGND VGND VPWR VPWR _02443_ sky130_fd_sc_hd__o221a_1
X_13639_ CPU.registerFile\[18\]\[22\] CPU.registerFile\[22\]\[22\] _07648_ VGND VGND
+ VPWR VPWR _08060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16358_ net2433 _07358_ _03829_ _03632_ VGND VGND VPWR VPWR _02441_ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15309_ _02797_ _02799_ _02801_ _02804_ _02807_ VGND VGND VPWR VPWR _02808_ sky130_fd_sc_hd__a221o_1
XFILLER_0_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16289_ _08408_ _03747_ _03762_ _08015_ VGND VGND VPWR VPWR _03763_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_117_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14910__993 clknet_1_1__leaf__02706_ VGND VGND VPWR VPWR net1025 sky130_fd_sc_hd__inv_2
X_18028_ net1201 _02308_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09801_ _05471_ VGND VGND VPWR VPWR _02524_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_130_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09732_ _04303_ _04698_ _04210_ _04300_ VGND VGND VPWR VPWR _05422_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_105_Left_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14527__648 clknet_1_0__leaf__02668_ VGND VGND VPWR VPWR net680 sky130_fd_sc_hd__inv_2
X_09663_ _05349_ _05355_ _04708_ VGND VGND VPWR VPWR _05356_ sky130_fd_sc_hd__o21ai_1
X_15065__1130 clknet_1_0__leaf__02723_ VGND VGND VPWR VPWR net1162 sky130_fd_sc_hd__inv_2
X_08614_ _04330_ _04256_ _04332_ _04333_ VGND VGND VPWR VPWR _04334_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09594_ net1274 CPU.instr\[2\] _04291_ _04830_ VGND VGND VPWR VPWR _05289_ sky130_fd_sc_hd__nand4_4
XFILLER_0_139_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08545_ CPU.aluIn1\[10\] _04263_ VGND VGND VPWR VPWR _04265_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08476_ CPU.instr\[3\] CPU.instr\[6\] CPU.instr\[4\] VGND VGND VPWR VPWR _04196_
+ sky130_fd_sc_hd__or3b_4
XFILLER_0_65_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_114_Left_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_150_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09028_ mapped_spi_ram.rcv_data\[3\] _04688_ _04709_ mapped_spi_flash.rcv_data\[3\]
+ VGND VGND VPWR VPWR _04744_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_14_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold260 CPU.cycles\[4\] VGND VGND VPWR VPWR net1501 sky130_fd_sc_hd__dlygate4sd3_1
X_14885__970 clknet_1_0__leaf__02704_ VGND VGND VPWR VPWR net1002 sky130_fd_sc_hd__inv_2
Xhold271 _02605_ VGND VGND VPWR VPWR net1512 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold282 CPU.rs2\[29\] VGND VGND VPWR VPWR net1523 sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 mapped_spi_ram.rcv_data\[15\] VGND VGND VPWR VPWR net1534 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Left_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_148_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12941_ _07281_ VGND VGND VPWR VPWR _07382_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_29_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15660_ _03065_ _03150_ _03151_ VGND VGND VPWR VPWR _03152_ sky130_fd_sc_hd__o21a_1
XANTENNA_100 _05381_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12872_ _07240_ VGND VGND VPWR VPWR _07314_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_158_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_111 _05425_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_122 _05528_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11823_ _06674_ VGND VGND VPWR VPWR _06675_ sky130_fd_sc_hd__buf_4
XANTENNA_133 _05551_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_144 _07253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15591_ CPU.registerFile\[12\]\[6\] _05049_ VGND VGND VPWR VPWR _03084_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_852 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_155 _07271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_166 _07325_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17330_ net519 _01618_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[26\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_177 _07476_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_885 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11754_ _05489_ _05775_ VGND VGND VPWR VPWR _06638_ sky130_fd_sc_hd__nand2_2
XANTENNA_188 _07841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_199 _07841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_132_Left_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10705_ _05511_ net2110 _06045_ VGND VGND VPWR VPWR _06046_ sky130_fd_sc_hd__mux2_1
X_17261_ net451 _01549_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[22\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_64_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14473_ clknet_1_1__leaf__02653_ VGND VGND VPWR VPWR _02663_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_81_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11685_ net1435 _06590_ _06595_ _06594_ VGND VGND VPWR VPWR _01713_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16212_ _02848_ _03683_ _03687_ _08410_ VGND VGND VPWR VPWR _03688_ sky130_fd_sc_hd__a211o_1
XFILLER_0_102_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13424_ CPU.registerFile\[8\]\[15\] CPU.registerFile\[12\]\[15\] _07318_ VGND VGND
+ VPWR VPWR _07852_ sky130_fd_sc_hd__mux2_1
X_17192_ clknet_leaf_25_clk _01480_ VGND VGND VPWR VPWR CPU.Iimm\[2\] sky130_fd_sc_hd__dfxtp_2
X_10636_ net1395 _05996_ _06002_ _05993_ VGND VGND VPWR VPWR _02172_ sky130_fd_sc_hd__o211a_1
Xclkload108 clknet_1_1__leaf__08357_ VGND VGND VPWR VPWR clkload108/Y sky130_fd_sc_hd__clkinvlp_4
X_16143_ CPU.registerFile\[1\]\[21\] _02939_ _03620_ _02894_ VGND VGND VPWR VPWR _03621_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13355_ _05284_ VGND VGND VPWR VPWR _07785_ sky130_fd_sc_hd__buf_6
XFILLER_0_122_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10567_ _05959_ _05952_ _05960_ net1507 VGND VGND VPWR VPWR _02199_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12306_ CPU.aluIn1\[3\] _06964_ _06859_ VGND VGND VPWR VPWR _06965_ sky130_fd_sc_hd__mux2_1
X_16074_ _03549_ _03553_ _03252_ VGND VGND VPWR VPWR _03554_ sky130_fd_sc_hd__a21o_1
X_13286_ CPU.registerFile\[5\]\[11\] _07373_ _07717_ _07368_ VGND VGND VPWR VPWR _07718_
+ sky130_fd_sc_hd__o211a_1
X_10498_ CPU.PC\[9\] _05867_ _05904_ _05905_ VGND VGND VPWR VPWR _05906_ sky130_fd_sc_hd__a22oi_2
X_12237_ _06912_ VGND VGND VPWR VPWR _01444_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_112_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12168_ CPU.aluWr _04681_ _06859_ VGND VGND VPWR VPWR _06860_ sky130_fd_sc_hd__a21oi_1
X_11119_ CPU.registerFile\[8\]\[19\] _05696_ _06263_ VGND VGND VPWR VPWR _06266_ sky130_fd_sc_hd__mux2_1
X_16976_ clknet_leaf_25_clk _01302_ VGND VGND VPWR VPWR CPU.mem_wdata\[7\] sky130_fd_sc_hd__dfxtp_2
X_12099_ _06821_ VGND VGND VPWR VPWR _01525_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14030__309 clknet_1_0__leaf__08362_ VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_88_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15927_ _08405_ _03409_ _03410_ VGND VGND VPWR VPWR _03411_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15858_ CPU.registerFile\[24\]\[13\] _03130_ _02790_ _03343_ VGND VGND VPWR VPWR
+ _03344_ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15789_ _02786_ _03274_ _03276_ _02794_ VGND VGND VPWR VPWR _03277_ sky130_fd_sc_hd__a211o_1
XFILLER_0_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17528_ net717 _01816_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17459_ net648 _01747_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_119_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09715_ _05404_ VGND VGND VPWR VPWR _05405_ sky130_fd_sc_hd__buf_6
X_09646_ mapped_spi_ram.rcv_data\[28\] net17 net1290 per_uart.rx_data\[4\] VGND VGND
+ VPWR VPWR _05339_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_143_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ _05272_ VGND VGND VPWR VPWR _05273_ sky130_fd_sc_hd__buf_4
XFILLER_0_78_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08528_ CPU.aluIn1\[19\] _04247_ VGND VGND VPWR VPWR _04248_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11470_ _05526_ net2477 _06444_ VGND VGND VPWR VPWR _06452_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10421_ net1347 _05841_ _05842_ net2538 _05844_ VGND VGND VPWR VPWR _02229_ sky130_fd_sc_hd__o221a_1
XFILLER_0_33_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13140_ _07256_ VGND VGND VPWR VPWR _07576_ sky130_fd_sc_hd__buf_4
XFILLER_0_61_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10352_ _05797_ VGND VGND VPWR VPWR _02252_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13071_ CPU.registerFile\[6\]\[5\] CPU.registerFile\[7\]\[5\] _07263_ VGND VGND VPWR
+ VPWR _07509_ sky130_fd_sc_hd__mux2_1
X_10283_ _05760_ VGND VGND VPWR VPWR _02299_ sky130_fd_sc_hd__clkbuf_1
X_12022_ _05426_ net1824 _06746_ VGND VGND VPWR VPWR _06780_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15113__1144 clknet_1_1__leaf__02724_ VGND VGND VPWR VPWR net1176 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16830_ _05816_ net20 _04130_ _04126_ net2100 VGND VGND VPWR VPWR _02612_ sky130_fd_sc_hd__a32o_1
X_16761_ _08436_ _08459_ _05063_ VGND VGND VPWR VPWR _04077_ sky130_fd_sc_hd__a21o_1
X_14248__420 clknet_1_1__leaf__08435_ VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__inv_2
X_15712_ CPU.registerFile\[1\]\[9\] _02867_ _03201_ _08405_ VGND VGND VPWR VPWR _03202_
+ sky130_fd_sc_hd__a22o_1
X_12924_ CPU.registerFile\[18\]\[2\] CPU.registerFile\[22\]\[2\] _07339_ VGND VGND
+ VPWR VPWR _07365_ sky130_fd_sc_hd__mux2_1
X_16692_ _04001_ _05298_ VGND VGND VPWR VPWR _04019_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_66_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12855_ CPU.registerFile\[28\]\[0\] CPU.registerFile\[24\]\[0\] _07297_ VGND VGND
+ VPWR VPWR _07298_ sky130_fd_sc_hd__mux2_1
X_15643_ CPU.registerFile\[29\]\[7\] _02800_ VGND VGND VPWR VPWR _03135_ sky130_fd_sc_hd__or2_1
X_11806_ _05273_ net2187 _06661_ VGND VGND VPWR VPWR _06666_ sky130_fd_sc_hd__mux2_1
X_15574_ _02831_ VGND VGND VPWR VPWR _03068_ sky130_fd_sc_hd__clkbuf_4
X_18362_ clknet_leaf_3_clk _02640_ VGND VGND VPWR VPWR per_uart.d_in_uart\[2\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12786_ _07228_ VGND VGND VPWR VPWR _07229_ sky130_fd_sc_hd__buf_2
XFILLER_0_28_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17313_ net502 _01601_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_16595__66 clknet_1_0__leaf__03970_ VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__inv_2
X_11737_ _06626_ VGND VGND VPWR VPWR _06627_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_56_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18293_ net126 _02573_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17244_ net434 _01532_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_12_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11668_ net1434 _06575_ _06585_ _06581_ VGND VGND VPWR VPWR _01720_ sky130_fd_sc_hd__o211a_1
XFILLER_0_142_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14556__674 clknet_1_1__leaf__02671_ VGND VGND VPWR VPWR net706 sky130_fd_sc_hd__inv_2
XFILLER_0_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13407_ CPU.registerFile\[18\]\[15\] CPU.registerFile\[22\]\[15\] _07233_ VGND VGND
+ VPWR VPWR _07835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17175_ clknet_leaf_24_clk _01463_ VGND VGND VPWR VPWR CPU.instr\[5\] sky130_fd_sc_hd__dfxtp_4
X_10619_ _05843_ VGND VGND VPWR VPWR _05993_ sky130_fd_sc_hd__buf_2
XFILLER_0_4_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11599_ _06508_ _06537_ VGND VGND VPWR VPWR _06538_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16126_ CPU.registerFile\[13\]\[21\] _03123_ VGND VGND VPWR VPWR _03604_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_114_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13338_ net1532 _07229_ _07768_ _07135_ VGND VGND VPWR VPWR _01307_ sky130_fd_sc_hd__o211a_1
X_16057_ CPU.registerFile\[21\]\[19\] CPU.registerFile\[23\]\[19\] _05441_ VGND VGND
+ VPWR VPWR _03537_ sky130_fd_sc_hd__mux2_1
X_13269_ _07411_ _07698_ _07701_ VGND VGND VPWR VPWR _07702_ sky130_fd_sc_hd__or3_1
Xclkbuf_1_1__f__02695_ clknet_0__02695_ VGND VGND VPWR VPWR clknet_1_1__leaf__02695_
+ sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__07222_ clknet_0__07222_ VGND VGND VPWR VPWR clknet_1_1__leaf__07222_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_138_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16959_ net254 _01285_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_09500_ _04264_ _04214_ _04219_ CPU.aluReg\[10\] _05198_ VGND VGND VPWR VPWR _05199_
+ sky130_fd_sc_hd__a221o_1
X_14721__822 clknet_1_0__leaf__02688_ VGND VGND VPWR VPWR net854 sky130_fd_sc_hd__inv_2
XFILLER_0_154_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09431_ _04710_ _05132_ _04636_ VGND VGND VPWR VPWR _05133_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09362_ _05067_ VGND VGND VPWR VPWR _02567_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14639__749 clknet_1_0__leaf__02679_ VGND VGND VPWR VPWR net781 sky130_fd_sc_hd__inv_2
XFILLER_0_47_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09293_ _04827_ _04828_ _04905_ VGND VGND VPWR VPWR _05002_ sky130_fd_sc_hd__and3_1
XANTENNA_11 _02852_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_22 _02940_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_33 _03100_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_44 _04696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_55 _04971_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_66 _05093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_77 _05170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_88 _05284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_99 _05380_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_113_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__03971_ clknet_0__03971_ VGND VGND VPWR VPWR clknet_1_0__leaf__03971_
+ sky130_fd_sc_hd__clkbuf_16
X_14384__519 clknet_1_1__leaf__02654_ VGND VGND VPWR VPWR net551 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_145_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap13 _06630_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_1
X_10970_ _06186_ VGND VGND VPWR VPWR _02023_ sky130_fd_sc_hd__clkbuf_1
Xmax_cap24 _04295_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__08360_ clknet_0__08360_ VGND VGND VPWR VPWR clknet_1_0__leaf__08360_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09629_ CPU.aluIn1\[5\] _04279_ _04211_ VGND VGND VPWR VPWR _05323_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_48_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12640_ _07144_ net1497 VGND VGND VPWR VPWR _00045_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12571_ CPU.registerFile\[4\]\[10\] _05208_ _07107_ VGND VGND VPWR VPWR _07109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_61_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11522_ mapped_spi_ram.snd_bitcount\[5\] mapped_spi_ram.snd_bitcount\[4\] mapped_spi_ram.snd_bitcount\[1\]
+ mapped_spi_ram.snd_bitcount\[0\] VGND VGND VPWR VPWR _06484_ sky130_fd_sc_hd__or4b_1
X_15290_ _05406_ VGND VGND VPWR VPWR _02789_ sky130_fd_sc_hd__buf_4
X_14850__939 clknet_1_0__leaf__02700_ VGND VGND VPWR VPWR net971 sky130_fd_sc_hd__inv_2
XFILLER_0_18_270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11453_ _05509_ net2233 _06433_ VGND VGND VPWR VPWR _06443_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10404_ _05832_ VGND VGND VPWR VPWR _02234_ sky130_fd_sc_hd__clkbuf_1
X_14172_ _08423_ VGND VGND VPWR VPWR _01486_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11384_ _06406_ VGND VGND VPWR VPWR _01829_ sky130_fd_sc_hd__clkbuf_1
X_13123_ CPU.registerFile\[29\]\[6\] _07556_ _07557_ CPU.registerFile\[25\]\[6\] _07559_
+ VGND VGND VPWR VPWR _07560_ sky130_fd_sc_hd__o221a_1
X_10335_ _05511_ net2111 _05788_ VGND VGND VPWR VPWR _05789_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ CPU.registerFile\[14\]\[4\] CPU.registerFile\[10\]\[4\] _07492_ VGND VGND
+ VPWR VPWR _07493_ sky130_fd_sc_hd__mux2_1
X_17931_ net1120 _02215_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[11\] sky130_fd_sc_hd__dfxtp_1
X_10266_ _05511_ net1757 _05751_ VGND VGND VPWR VPWR _05752_ sky130_fd_sc_hd__mux2_1
X_12005_ _06771_ VGND VGND VPWR VPWR _01570_ sky130_fd_sc_hd__clkbuf_1
X_17862_ net1051 _02146_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10197_ _05707_ VGND VGND VPWR VPWR _02332_ sky130_fd_sc_hd__clkbuf_1
X_16813_ _07177_ _08355_ VGND VGND VPWR VPWR _04118_ sky130_fd_sc_hd__nor2_1
X_17793_ net982 _02077_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16744_ _04052_ _05127_ _04006_ VGND VGND VPWR VPWR _04063_ sky130_fd_sc_hd__or3b_1
X_12907_ _04971_ VGND VGND VPWR VPWR _07349_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_17_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16675_ _03991_ net1539 VGND VGND VPWR VPWR _04004_ sky130_fd_sc_hd__nand2_1
X_13887_ CPU.registerFile\[16\]\[30\] CPU.registerFile\[20\]\[30\] _07314_ VGND VGND
+ VPWR VPWR _08300_ sky130_fd_sc_hd__mux2_1
X_15626_ _02772_ VGND VGND VPWR VPWR _03118_ sky130_fd_sc_hd__clkbuf_2
X_12838_ _07235_ VGND VGND VPWR VPWR _07281_ sky130_fd_sc_hd__buf_4
XFILLER_0_118_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18345_ clknet_leaf_1_clk _02625_ VGND VGND VPWR VPWR per_uart.uart0.rx_busy sky130_fd_sc_hd__dfxtp_1
X_15557_ CPU.registerFile\[27\]\[5\] CPU.registerFile\[31\]\[5\] _03050_ VGND VGND
+ VPWR VPWR _03051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15488_ _02979_ _02981_ _02983_ _02945_ VGND VGND VPWR VPWR _02984_ sky130_fd_sc_hd__o22a_1
X_18276_ net109 _02556_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__03965_ _03965_ VGND VGND VPWR VPWR clknet_0__03965_ sky130_fd_sc_hd__clkbuf_16
X_17227_ net417 _01515_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_96_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17158_ net382 _01446_ VGND VGND VPWR VPWR CPU.aluReg\[22\] sky130_fd_sc_hd__dfxtp_1
Xhold804 CPU.registerFile\[30\]\[13\] VGND VGND VPWR VPWR net2045 sky130_fd_sc_hd__dlygate4sd3_1
Xhold815 CPU.registerFile\[2\]\[2\] VGND VGND VPWR VPWR net2056 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold826 CPU.registerFile\[29\]\[29\] VGND VGND VPWR VPWR net2067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold837 CPU.registerFile\[23\]\[31\] VGND VGND VPWR VPWR net2078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold848 CPU.registerFile\[15\]\[20\] VGND VGND VPWR VPWR net2089 sky130_fd_sc_hd__dlygate4sd3_1
X_16109_ _03583_ _03587_ _02784_ VGND VGND VPWR VPWR _03588_ sky130_fd_sc_hd__a21o_1
X_09980_ _05535_ net2403 _05581_ VGND VGND VPWR VPWR _05583_ sky130_fd_sc_hd__mux2_1
X_17089_ net347 _01411_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[19\] sky130_fd_sc_hd__dfxtp_1
Xhold859 per_uart.uart0.tx_bitcount\[1\] VGND VGND VPWR VPWR net2100 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__02747_ clknet_0__02747_ VGND VGND VPWR VPWR clknet_1_1__leaf__02747_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08931_ _04625_ _04622_ _04650_ _04649_ VGND VGND VPWR VPWR _04651_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__02678_ clknet_0__02678_ VGND VGND VPWR VPWR clknet_1_1__leaf__02678_
+ sky130_fd_sc_hd__clkbuf_16
X_08862_ _04581_ CPU.aluIn1\[23\] VGND VGND VPWR VPWR _04582_ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_127_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08793_ CPU.aluIn1\[8\] CPU.Bimm\[8\] VGND VGND VPWR VPWR _04513_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_127_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09414_ _04258_ _04699_ _04808_ CPU.aluReg\[14\] _05116_ VGND VGND VPWR VPWR _05117_
+ sky130_fd_sc_hd__a221o_1
X_16559__33 clknet_1_0__leaf__03967_ VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__inv_2
XFILLER_0_48_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09345_ _04504_ _05050_ _04777_ VGND VGND VPWR VPWR _05051_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15112__1143 clknet_1_1__leaf__02724_ VGND VGND VPWR VPWR net1175 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_43_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09276_ mapped_spi_ram.rcv_data\[12\] _04688_ _04690_ mapped_spi_flash.rcv_data\[12\]
+ VGND VGND VPWR VPWR _04985_ sky130_fd_sc_hd__a22oi_4
X_16574__47 clknet_1_1__leaf__03968_ VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__inv_2
XFILLER_0_74_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10120_ net2361 _05230_ _05655_ VGND VGND VPWR VPWR _05658_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10051_ net2239 _05230_ _05618_ VGND VGND VPWR VPWR _05621_ sky130_fd_sc_hd__mux2_1
X_13810_ CPU.registerFile\[30\]\[27\] CPU.registerFile\[26\]\[27\] _07292_ VGND VGND
+ VPWR VPWR _08226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13741_ CPU.registerFile\[18\]\[25\] CPU.registerFile\[22\]\[25\] _05283_ VGND VGND
+ VPWR VPWR _08159_ sky130_fd_sc_hd__mux2_1
X_10953_ net1673 _05735_ _06142_ VGND VGND VPWR VPWR _06177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16460_ CPU.registerFile\[5\]\[31\] CPU.registerFile\[4\]\[31\] _05092_ VGND VGND
+ VPWR VPWR _03928_ sky130_fd_sc_hd__mux2_1
X_13672_ CPU.registerFile\[18\]\[23\] CPU.registerFile\[22\]\[23\] _07648_ VGND VGND
+ VPWR VPWR _08092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_816 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10884_ net1622 _05735_ _06105_ VGND VGND VPWR VPWR _06140_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_155_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15411_ CPU.registerFile\[8\]\[2\] CPU.registerFile\[12\]\[2\] _08403_ VGND VGND
+ VPWR VPWR _02908_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__02698_ clknet_0__02698_ VGND VGND VPWR VPWR clknet_1_0__leaf__02698_
+ sky130_fd_sc_hd__clkbuf_16
X_12623_ net1328 net1492 VGND VGND VPWR VPWR _00026_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_158_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16391_ _08407_ _03838_ _03847_ _03861_ _07424_ VGND VGND VPWR VPWR _03862_ sky130_fd_sc_hd__a311o_1
XFILLER_0_155_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__07225_ clknet_0__07225_ VGND VGND VPWR VPWR clknet_1_0__leaf__07225_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_158_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_23_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_8
X_18130_ net193 _02410_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_15342_ _02827_ _02839_ _02840_ VGND VGND VPWR VPWR _02841_ sky130_fd_sc_hd__o21ai_1
X_12554_ net2044 _05045_ _07096_ VGND VGND VPWR VPWR _07100_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11505_ mapped_spi_ram.state\[2\] mapped_spi_ram.state\[0\] VGND VGND VPWR VPWR _06472_
+ sky130_fd_sc_hd__nor2_1
X_18061_ net1234 _02341_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_15273_ _05048_ VGND VGND VPWR VPWR _02772_ sky130_fd_sc_hd__buf_4
X_12485_ _07063_ VGND VGND VPWR VPWR _01347_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17012_ net270 _01334_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_78_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14224_ clknet_1_0__leaf__08363_ VGND VGND VPWR VPWR _08432_ sky130_fd_sc_hd__buf_1
XFILLER_0_62_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11436_ _06434_ VGND VGND VPWR VPWR _01805_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__02701_ _02701_ VGND VGND VPWR VPWR clknet_0__02701_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_123_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14155_ _08414_ VGND VGND VPWR VPWR _01478_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11367_ _05487_ net1868 _06397_ VGND VGND VPWR VPWR _06398_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13106_ CPU.registerFile\[6\]\[6\] _05337_ VGND VGND VPWR VPWR _07543_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10318_ _05495_ net2238 _05777_ VGND VGND VPWR VPWR _05780_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11298_ _05487_ net2078 _06360_ VGND VGND VPWR VPWR _06361_ sky130_fd_sc_hd__mux2_1
X_14668__775 clknet_1_1__leaf__02682_ VGND VGND VPWR VPWR net807 sky130_fd_sc_hd__inv_2
X_13037_ _07352_ VGND VGND VPWR VPWR _07476_ sky130_fd_sc_hd__buf_8
X_17914_ net1103 _02198_ VGND VGND VPWR VPWR mapped_spi_flash.snd_bitcount\[0\] sky130_fd_sc_hd__dfxtp_1
X_10249_ _05495_ net2170 _05740_ VGND VGND VPWR VPWR _05743_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17845_ net1034 _02129_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_109_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17776_ net965 _02060_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16727_ _04044_ _04048_ _04015_ VGND VGND VPWR VPWR _02591_ sky130_fd_sc_hd__a21oi_1
X_13939_ _07330_ _08350_ VGND VGND VPWR VPWR _08351_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_122_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15609_ CPU.registerFile\[1\]\[6\] _02814_ _03101_ _02816_ VGND VGND VPWR VPWR _03102_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_158_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_14_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_84_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14833__923 clknet_1_1__leaf__02699_ VGND VGND VPWR VPWR net955 sky130_fd_sc_hd__inv_2
XFILLER_0_56_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09130_ CPU.Jimm\[16\] _04829_ _04831_ VGND VGND VPWR VPWR _04842_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18328_ clknet_leaf_5_clk _02608_ VGND VGND VPWR VPWR per_uart.uart0.tx_count16\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09061_ CPU.Bimm\[5\] _04498_ _04503_ CPU.cycles\[25\] VGND VGND VPWR VPWR _04775_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_100_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18259_ net100 _02539_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold601 CPU.registerFile\[1\]\[29\] VGND VGND VPWR VPWR net1842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold612 CPU.registerFile\[15\]\[24\] VGND VGND VPWR VPWR net1853 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold623 CPU.registerFile\[14\]\[13\] VGND VGND VPWR VPWR net1864 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold634 CPU.registerFile\[26\]\[19\] VGND VGND VPWR VPWR net1875 sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 CPU.registerFile\[16\]\[5\] VGND VGND VPWR VPWR net1886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold656 CPU.registerFile\[9\]\[24\] VGND VGND VPWR VPWR net1897 sky130_fd_sc_hd__dlygate4sd3_1
Xhold667 CPU.registerFile\[29\]\[15\] VGND VGND VPWR VPWR net1908 sky130_fd_sc_hd__dlygate4sd3_1
X_09963_ _05518_ net1612 _05570_ VGND VGND VPWR VPWR _05574_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold678 CPU.registerFile\[29\]\[0\] VGND VGND VPWR VPWR net1919 sky130_fd_sc_hd__dlygate4sd3_1
Xhold689 mapped_spi_ram.cmd_addr\[0\] VGND VGND VPWR VPWR net1930 sky130_fd_sc_hd__dlygate4sd3_1
X_08914_ _04520_ _04632_ VGND VGND VPWR VPWR _04634_ sky130_fd_sc_hd__nand2_1
X_09894_ _05530_ net2042 _05512_ VGND VGND VPWR VPWR _05531_ sky130_fd_sc_hd__mux2_1
Xhold1301 mapped_spi_ram.rcv_bitcount\[1\] VGND VGND VPWR VPWR net2542 sky130_fd_sc_hd__dlygate4sd3_1
X_08845_ CPU.aluIn1\[19\] _04495_ VGND VGND VPWR VPWR _04565_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_0__07219_ _07219_ VGND VGND VPWR VPWR clknet_0__07219_ sky130_fd_sc_hd__clkbuf_16
X_08776_ _04495_ VGND VGND VPWR VPWR _04496_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_0_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09328_ _04445_ _05034_ VGND VGND VPWR VPWR _05035_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_105_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09259_ CPU.cycles\[21\] _04503_ _04968_ _04773_ VGND VGND VPWR VPWR _04969_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_153_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12270_ CPU.aluReg\[12\] _06937_ _06924_ VGND VGND VPWR VPWR _06938_ sky130_fd_sc_hd__mux2_1
X_11221_ _06319_ VGND VGND VPWR VPWR _01905_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11152_ CPU.registerFile\[8\]\[3\] _05729_ _06274_ VGND VGND VPWR VPWR _06283_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10103_ net2267 _05066_ _05644_ VGND VGND VPWR VPWR _05649_ sky130_fd_sc_hd__mux2_1
X_11083_ net2217 _05729_ _06237_ VGND VGND VPWR VPWR _06246_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15960_ _02911_ _03440_ _03442_ _03245_ VGND VGND VPWR VPWR _03443_ sky130_fd_sc_hd__a211o_1
X_10034_ net2386 _05066_ _05607_ VGND VGND VPWR VPWR _05612_ sky130_fd_sc_hd__mux2_1
X_15891_ CPU.registerFile\[28\]\[14\] _03064_ VGND VGND VPWR VPWR _03376_ sky130_fd_sc_hd__or2_1
X_17630_ net819 _01918_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_15217__128 clknet_1_0__leaf__02752_ VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__inv_2
X_17561_ net750 _01849_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_14773_ clknet_1_0__leaf__02686_ VGND VGND VPWR VPWR _02693_ sky130_fd_sc_hd__buf_1
X_11985_ _05027_ net2048 _06758_ VGND VGND VPWR VPWR _06761_ sky130_fd_sc_hd__mux2_1
X_10936_ _06168_ VGND VGND VPWR VPWR _02039_ sky130_fd_sc_hd__clkbuf_1
X_13724_ CPU.registerFile\[28\]\[25\] CPU.registerFile\[24\]\[25\] _04938_ VGND VGND
+ VPWR VPWR _08142_ sky130_fd_sc_hd__mux2_1
X_17492_ net681 _01780_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_27_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16443_ CPU.registerFile\[28\]\[30\] CPU.registerFile\[24\]\[30\] _02881_ VGND VGND
+ VPWR VPWR _03912_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10867_ _06131_ VGND VGND VPWR VPWR _02071_ sky130_fd_sc_hd__clkbuf_1
X_13655_ CPU.registerFile\[29\]\[22\] _07347_ _07348_ CPU.registerFile\[25\]\[22\]
+ _08075_ VGND VGND VPWR VPWR _08076_ sky130_fd_sc_hd__o221a_1
X_16538__14 clknet_1_0__leaf__03965_ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__inv_2
XFILLER_0_128_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_144_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12606_ _07125_ _05970_ _06016_ _05942_ VGND VGND VPWR VPWR _00007_ sky130_fd_sc_hd__o31a_1
XFILLER_0_54_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16374_ CPU.registerFile\[25\]\[28\] _03280_ _02940_ VGND VGND VPWR VPWR _03845_
+ sky130_fd_sc_hd__o21a_1
X_13586_ CPU.registerFile\[31\]\[20\] _07556_ _07557_ CPU.registerFile\[27\]\[20\]
+ _08008_ VGND VGND VPWR VPWR _08009_ sky130_fd_sc_hd__o221a_1
XFILLER_0_143_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10798_ _05537_ net1804 _06092_ VGND VGND VPWR VPWR _06095_ sky130_fd_sc_hd__mux2_1
X_18113_ net176 _02393_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15325_ _02818_ _02820_ _02823_ VGND VGND VPWR VPWR _02824_ sky130_fd_sc_hd__a21o_1
X_12537_ net2483 _04761_ _07085_ VGND VGND VPWR VPWR _07091_ sky130_fd_sc_hd__mux2_1
X_16553__28 clknet_1_0__leaf__03966_ VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__inv_2
XFILLER_0_81_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18044_ net1217 _02324_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_12468_ _07054_ VGND VGND VPWR VPWR _01355_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11419_ _05543_ net2051 _06419_ VGND VGND VPWR VPWR _06425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12399_ _04748_ net2277 _07013_ VGND VGND VPWR VPWR _07018_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14138_ CPU.Jimm\[16\] _08401_ _08387_ VGND VGND VPWR VPWR _08402_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_3_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_8
X_08630_ _04236_ _04349_ VGND VGND VPWR VPWR _04350_ sky130_fd_sc_hd__nor2_1
X_17828_ net1017 _02112_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08561_ CPU.aluIn1\[5\] _04279_ VGND VGND VPWR VPWR _04281_ sky130_fd_sc_hd__or2_1
X_17759_ net948 _02043_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_703 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08492_ CPU.aluIn1\[31\] _04207_ _04211_ VGND VGND VPWR VPWR _04212_ sky130_fd_sc_hd__o21a_1
XFILLER_0_65_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14421__552 clknet_1_1__leaf__02658_ VGND VGND VPWR VPWR net584 sky130_fd_sc_hd__inv_2
XFILLER_0_18_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_135_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09113_ _04823_ _04824_ VGND VGND VPWR VPWR _04825_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09044_ _04216_ _04758_ _04655_ VGND VGND VPWR VPWR _04759_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_115_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14339__479 clknet_1_1__leaf__08466_ VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__inv_2
XFILLER_0_5_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold420 CPU.registerFile\[28\]\[20\] VGND VGND VPWR VPWR net1661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 CPU.registerFile\[6\]\[21\] VGND VGND VPWR VPWR net1672 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold442 CPU.registerFile\[30\]\[3\] VGND VGND VPWR VPWR net1683 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold453 CPU.registerFile\[18\]\[2\] VGND VGND VPWR VPWR net1694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 CPU.registerFile\[19\]\[10\] VGND VGND VPWR VPWR net1705 sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 CPU.registerFile\[15\]\[0\] VGND VGND VPWR VPWR net1716 sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 CPU.registerFile\[5\]\[24\] VGND VGND VPWR VPWR net1727 sky130_fd_sc_hd__dlygate4sd3_1
Xhold497 CPU.registerFile\[28\]\[17\] VGND VGND VPWR VPWR net1738 sky130_fd_sc_hd__dlygate4sd3_1
X_09946_ _05501_ net1651 _05559_ VGND VGND VPWR VPWR _05565_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_5_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ _05519_ VGND VGND VPWR VPWR _02496_ sky130_fd_sc_hd__clkbuf_1
Xhold1120 CPU.registerFile\[18\]\[9\] VGND VGND VPWR VPWR net2361 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1131 CPU.registerFile\[27\]\[17\] VGND VGND VPWR VPWR net2372 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1142 CPU.registerFile\[18\]\[16\] VGND VGND VPWR VPWR net2383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1153 CPU.registerFile\[15\]\[21\] VGND VGND VPWR VPWR net2394 sky130_fd_sc_hd__dlygate4sd3_1
X_08828_ _04511_ _04547_ VGND VGND VPWR VPWR _04548_ sky130_fd_sc_hd__and2_4
Xhold1164 CPU.registerFile\[12\]\[15\] VGND VGND VPWR VPWR net2405 sky130_fd_sc_hd__dlygate4sd3_1
X_14805__899 clknet_1_0__leaf__02695_ VGND VGND VPWR VPWR net931 sky130_fd_sc_hd__inv_2
Xhold1175 CPU.registerFile\[11\]\[22\] VGND VGND VPWR VPWR net2416 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1186 CPU.PC\[10\] VGND VGND VPWR VPWR net2427 sky130_fd_sc_hd__dlygate4sd3_1
X_08759_ CPU.aluIn1\[30\] VGND VGND VPWR VPWR _04479_ sky130_fd_sc_hd__inv_2
Xhold1197 CPU.registerFile\[15\]\[27\] VGND VGND VPWR VPWR net2438 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_304 _07404_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_315 _07914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14049__325 clknet_1_0__leaf__08365_ VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__inv_2
X_14504__627 clknet_1_1__leaf__02666_ VGND VGND VPWR VPWR net659 sky130_fd_sc_hd__inv_2
XANTENNA_326 _07930_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_337 _02895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11770_ _04798_ net1954 _06639_ VGND VGND VPWR VPWR _06647_ sky130_fd_sc_hd__mux2_1
XANTENNA_348 _05338_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_359 _07268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14242__415 clknet_1_0__leaf__08434_ VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__inv_2
X_10721_ _05528_ net1601 _06045_ VGND VGND VPWR VPWR _06054_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13440_ CPU.registerFile\[16\]\[16\] CPU.registerFile\[20\]\[16\] _07258_ VGND VGND
+ VPWR VPWR _07867_ sky130_fd_sc_hd__mux2_1
X_10652_ _06010_ _06011_ VGND VGND VPWR VPWR _06012_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13371_ net1526 _07229_ _07800_ _07135_ VGND VGND VPWR VPWR _01308_ sky130_fd_sc_hd__o211a_1
X_10583_ net1453 _05970_ VGND VGND VPWR VPWR _05973_ sky130_fd_sc_hd__or2_1
X_15110_ _05843_ per_uart.uart0.enable16_counter\[15\] _07193_ VGND VGND VPWR VPWR
+ _02742_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12322_ _06976_ VGND VGND VPWR VPWR _06977_ sky130_fd_sc_hd__buf_4
X_16090_ CPU.registerFile\[2\]\[20\] _03227_ _03228_ CPU.registerFile\[3\]\[20\] _03568_
+ VGND VGND VPWR VPWR _03569_ sky130_fd_sc_hd__a221o_1
XFILLER_0_121_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15041_ clknet_1_1__leaf__07222_ VGND VGND VPWR VPWR _02720_ sky130_fd_sc_hd__buf_1
XFILLER_0_121_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12253_ CPU.aluReg\[16\] _06923_ _06924_ VGND VGND VPWR VPWR _06925_ sky130_fd_sc_hd__mux2_1
X_14550__669 clknet_1_1__leaf__02670_ VGND VGND VPWR VPWR net701 sky130_fd_sc_hd__inv_2
X_11204_ _05532_ net2183 _06310_ VGND VGND VPWR VPWR _06311_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12184_ _06870_ VGND VGND VPWR VPWR _06871_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_71_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11135_ _06251_ VGND VGND VPWR VPWR _06274_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16992_ clknet_leaf_28_clk _01318_ VGND VGND VPWR VPWR CPU.rs2\[23\] sky130_fd_sc_hd__dfxtp_1
X_11066_ _06214_ VGND VGND VPWR VPWR _06237_ sky130_fd_sc_hd__clkbuf_4
X_15943_ CPU.registerFile\[16\]\[15\] CPU.registerFile\[18\]\[15\] _03032_ VGND VGND
+ VPWR VPWR _03427_ sky130_fd_sc_hd__mux2_1
X_10017_ net2195 _04780_ _05596_ VGND VGND VPWR VPWR _05603_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15874_ CPU.registerFile\[22\]\[13\] CPU.registerFile\[23\]\[13\] _02828_ VGND VGND
+ VPWR VPWR _03360_ sky130_fd_sc_hd__mux2_1
X_17613_ net802 _01901_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17544_ net733 _01832_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_102_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11968_ _04748_ net2193 _06747_ VGND VGND VPWR VPWR _06752_ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13707_ _07646_ _08115_ _08118_ _08125_ VGND VGND VPWR VPWR _08126_ sky130_fd_sc_hd__a31o_1
X_10919_ _06159_ VGND VGND VPWR VPWR _02047_ sky130_fd_sc_hd__clkbuf_1
X_17475_ net664 _01763_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[30\] sky130_fd_sc_hd__dfxtp_1
X_11899_ _06715_ VGND VGND VPWR VPWR _01620_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16426_ _02757_ _03886_ _03895_ _07308_ VGND VGND VPWR VPWR _03896_ sky130_fd_sc_hd__a31o_1
XFILLER_0_39_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13638_ _07273_ _08057_ _08058_ VGND VGND VPWR VPWR _08059_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16357_ _02879_ _03810_ _03828_ _02846_ VGND VGND VPWR VPWR _03829_ sky130_fd_sc_hd__a211o_1
X_13569_ CPU.registerFile\[1\]\[20\] _07387_ _07991_ _07379_ VGND VGND VPWR VPWR _07992_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_70_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15308_ _02806_ VGND VGND VPWR VPWR _02807_ sky130_fd_sc_hd__buf_4
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16288_ _03755_ _03761_ _02844_ VGND VGND VPWR VPWR _03762_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_117_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18027_ net1200 _02307_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09800_ net2242 _05130_ _05463_ VGND VGND VPWR VPWR _05471_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_130_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09731_ _05415_ _04701_ VGND VGND VPWR VPWR _05421_ sky130_fd_sc_hd__nor2_1
X_09662_ _04419_ _04806_ _05354_ _04768_ VGND VGND VPWR VPWR _05355_ sky130_fd_sc_hd__a2bb2o_1
X_08613_ CPU.aluIn1\[16\] _04254_ VGND VGND VPWR VPWR _04333_ sky130_fd_sc_hd__xnor2_1
X_09593_ _04500_ VGND VGND VPWR VPWR _05288_ sky130_fd_sc_hd__buf_2
XFILLER_0_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08544_ CPU.aluIn1\[10\] _04263_ VGND VGND VPWR VPWR _04264_ sky130_fd_sc_hd__and2_1
X_08475_ _04195_ VGND VGND VPWR VPWR _02646_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_476 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15246__154 clknet_1_1__leaf__02755_ VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__inv_2
X_09027_ _04359_ _04489_ _04739_ _04742_ VGND VGND VPWR VPWR _04743_ sky130_fd_sc_hd__a211o_1
XFILLER_0_14_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold250 CPU.cycles\[22\] VGND VGND VPWR VPWR net1491 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold261 CPU.cycles\[25\] VGND VGND VPWR VPWR net1502 sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 CPU.state\[1\] VGND VGND VPWR VPWR net1513 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold283 CPU.cycles\[15\] VGND VGND VPWR VPWR net1524 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 CPU.rs2\[21\] VGND VGND VPWR VPWR net1535 sky130_fd_sc_hd__dlygate4sd3_1
X_09929_ _05554_ VGND VGND VPWR VPWR _02479_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_130_Right_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_148_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12940_ _07360_ _07367_ _07378_ _07380_ VGND VGND VPWR VPWR _07381_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ CPU.registerFile\[6\]\[1\] CPU.registerFile\[7\]\[1\] _07263_ VGND VGND VPWR
+ VPWR _07313_ sky130_fd_sc_hd__mux2_1
XANTENNA_101 _05381_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_112 _05425_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_123 _05530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11822_ _05631_ _06250_ VGND VGND VPWR VPWR _06674_ sky130_fd_sc_hd__nor2_2
XANTENNA_134 _05694_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15590_ CPU.registerFile\[14\]\[6\] CPU.registerFile\[10\]\[6\] _03082_ VGND VGND
+ VPWR VPWR _03083_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_145 _07253_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_156 _07271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_167 _07326_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_139_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_178 _07480_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11753_ net1505 _06627_ _06635_ VGND VGND VPWR VPWR _01688_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_189 _07841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10704_ _06033_ VGND VGND VPWR VPWR _06045_ sky130_fd_sc_hd__buf_4
X_17260_ net450 _01548_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11684_ mapped_spi_ram.rcv_data\[18\] _06588_ VGND VGND VPWR VPWR _06595_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16211_ _02856_ _03684_ _03686_ _03019_ VGND VGND VPWR VPWR _03687_ sky130_fd_sc_hd__o211a_1
X_13423_ _07818_ _07849_ _07850_ VGND VGND VPWR VPWR _07851_ sky130_fd_sc_hd__o21a_1
X_10635_ mapped_spi_flash.rcv_data\[6\] _05994_ VGND VGND VPWR VPWR _06002_ sky130_fd_sc_hd__or2_1
X_17191_ clknet_leaf_25_clk _01479_ VGND VGND VPWR VPWR CPU.Iimm\[1\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_52_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload109 clknet_1_0__leaf__08356_ VGND VGND VPWR VPWR clkload109/Y sky130_fd_sc_hd__clkinvlp_4
X_13354_ _07777_ _07783_ _04814_ VGND VGND VPWR VPWR _07784_ sky130_fd_sc_hd__mux2_1
X_16142_ CPU.registerFile\[5\]\[21\] CPU.registerFile\[4\]\[21\] _03146_ VGND VGND
+ VPWR VPWR _03620_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10566_ _05850_ mapped_spi_flash.snd_bitcount\[0\] _05950_ VGND VGND VPWR VPWR _05960_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12305_ CPU.aluReg\[4\] CPU.aluReg\[2\] _06939_ VGND VGND VPWR VPWR _06964_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13285_ CPU.registerFile\[4\]\[11\] _07388_ VGND VGND VPWR VPWR _07717_ sky130_fd_sc_hd__or2_1
X_16073_ _02924_ _03550_ _03551_ _03552_ _02782_ VGND VGND VPWR VPWR _03553_ sky130_fd_sc_hd__a221o_1
X_10497_ _05903_ _04544_ _04543_ _04590_ VGND VGND VPWR VPWR _05905_ sky130_fd_sc_hd__o31a_1
XFILLER_0_32_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12236_ net2470 _06911_ _06891_ VGND VGND VPWR VPWR _06912_ sky130_fd_sc_hd__mux2_1
X_12167_ _06858_ VGND VGND VPWR VPWR _06859_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_112_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11118_ _06265_ VGND VGND VPWR VPWR _01954_ sky130_fd_sc_hd__clkbuf_1
X_16975_ clknet_leaf_22_clk _01301_ VGND VGND VPWR VPWR CPU.mem_wdata\[6\] sky130_fd_sc_hd__dfxtp_2
X_12098_ _04696_ net2387 _06819_ VGND VGND VPWR VPWR _06821_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15926_ CPU.registerFile\[2\]\[15\] _02872_ _02873_ CPU.registerFile\[3\]\[15\] _02875_
+ VGND VGND VPWR VPWR _03410_ sky130_fd_sc_hd__a221o_1
X_11049_ _06228_ VGND VGND VPWR VPWR _01986_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15857_ CPU.registerFile\[28\]\[13\] _03064_ VGND VGND VPWR VPWR _03343_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15788_ CPU.registerFile\[24\]\[11\] _03130_ _02790_ _03275_ VGND VGND VPWR VPWR
+ _03276_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17527_ net716 _01815_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17458_ net647 _01746_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_119_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16409_ CPU.registerFile\[14\]\[29\] _02889_ VGND VGND VPWR VPWR _03879_ sky130_fd_sc_hd__or2_1
XFILLER_0_144_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17389_ net578 _01677_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_99_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14078__351 clknet_1_0__leaf__08368_ VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__inv_2
XFILLER_0_2_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14533__653 clknet_1_1__leaf__02669_ VGND VGND VPWR VPWR net685 sky130_fd_sc_hd__inv_2
XFILLER_0_11_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09714_ mapped_spi_ram.rcv_data\[9\] net18 _04690_ mapped_spi_flash.rcv_data\[9\]
+ VGND VGND VPWR VPWR _05404_ sky130_fd_sc_hd__a22o_1
X_14189__368 clknet_1_0__leaf__08428_ VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__inv_2
X_09645_ _05337_ VGND VGND VPWR VPWR _05338_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_117_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09576_ CPU.cycles\[7\] _04687_ _05271_ VGND VGND VPWR VPWR _05272_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_143_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ CPU.rs2\[19\] _04200_ _04205_ VGND VGND VPWR VPWR _04247_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14616__728 clknet_1_1__leaf__02677_ VGND VGND VPWR VPWR net760 sky130_fd_sc_hd__inv_2
XFILLER_0_18_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10420_ _05843_ VGND VGND VPWR VPWR _05844_ sky130_fd_sc_hd__buf_4
XFILLER_0_61_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10351_ _05528_ net2060 _05788_ VGND VGND VPWR VPWR _05797_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13070_ CPU.registerFile\[2\]\[5\] CPU.registerFile\[3\]\[5\] _07311_ VGND VGND VPWR
+ VPWR _07508_ sky130_fd_sc_hd__mux2_1
X_10282_ _05528_ net1931 _05751_ VGND VGND VPWR VPWR _05760_ sky130_fd_sc_hd__mux2_1
X_12021_ _06779_ VGND VGND VPWR VPWR _01562_ sky130_fd_sc_hd__clkbuf_1
X_16760_ _03990_ CPU.PC\[17\] VGND VGND VPWR VPWR _04076_ sky130_fd_sc_hd__and2_1
X_15711_ CPU.registerFile\[5\]\[9\] CPU.registerFile\[4\]\[9\] _02806_ VGND VGND VPWR
+ VPWR _03201_ sky130_fd_sc_hd__mux2_1
X_12923_ _07245_ VGND VGND VPWR VPWR _07364_ sky130_fd_sc_hd__buf_2
X_16691_ _05288_ _05292_ _08454_ VGND VGND VPWR VPWR _04018_ sky130_fd_sc_hd__and3_1
XFILLER_0_158_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15642_ CPU.registerFile\[27\]\[7\] CPU.registerFile\[31\]\[7\] _03050_ VGND VGND
+ VPWR VPWR _03134_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ _04937_ VGND VGND VPWR VPWR _07297_ sky130_fd_sc_hd__buf_4
X_11805_ _06665_ VGND VGND VPWR VPWR _01664_ sky130_fd_sc_hd__clkbuf_1
X_18361_ clknet_leaf_3_clk _02639_ VGND VGND VPWR VPWR per_uart.d_in_uart\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15573_ CPU.registerFile\[20\]\[5\] CPU.registerFile\[21\]\[5\] _03066_ VGND VGND
+ VPWR VPWR _03067_ sky130_fd_sc_hd__mux2_1
X_12785_ _07227_ VGND VGND VPWR VPWR _07228_ sky130_fd_sc_hd__buf_2
XFILLER_0_84_823 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17312_ net501 _01600_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18292_ net125 _02572_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_11736_ _06471_ _06625_ _00008_ VGND VGND VPWR VPWR _06626_ sky130_fd_sc_hd__or3_1
XFILLER_0_154_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17243_ net433 _01531_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_12_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11667_ net1322 _06577_ VGND VGND VPWR VPWR _06585_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13406_ net1548 _07229_ _07834_ _07135_ VGND VGND VPWR VPWR _01309_ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17174_ clknet_leaf_24_clk _01462_ VGND VGND VPWR VPWR CPU.instr\[4\] sky130_fd_sc_hd__dfxtp_1
X_10618_ mapped_spi_flash.rcv_data\[13\] _05981_ VGND VGND VPWR VPWR _05992_ sky130_fd_sc_hd__or2_1
X_11598_ _04639_ net1350 _06493_ VGND VGND VPWR VPWR _06537_ sky130_fd_sc_hd__mux2_1
X_16125_ CPU.registerFile\[15\]\[21\] CPU.registerFile\[11\]\[21\] _02906_ VGND VGND
+ VPWR VPWR _03603_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13337_ _07230_ _07752_ _07767_ _07309_ VGND VGND VPWR VPWR _07768_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_114_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10549_ mapped_spi_flash.snd_bitcount\[5\] _05945_ VGND VGND VPWR VPWR _05947_ sky130_fd_sc_hd__or2_1
X_16056_ _03532_ _03535_ _02858_ VGND VGND VPWR VPWR _03536_ sky130_fd_sc_hd__mux2_2
XFILLER_0_11_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13268_ _07475_ _07699_ _07700_ VGND VGND VPWR VPWR _07701_ sky130_fd_sc_hd__o21a_1
Xclkbuf_1_1__f__02694_ clknet_0__02694_ VGND VGND VPWR VPWR clknet_1_1__leaf__02694_
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f__07221_ clknet_0__07221_ VGND VGND VPWR VPWR clknet_1_1__leaf__07221_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_94_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12219_ CPU.aluReg\[24\] _06898_ _06891_ VGND VGND VPWR VPWR _06899_ sky130_fd_sc_hd__mux2_1
X_13199_ _07475_ _07632_ _07633_ VGND VGND VPWR VPWR _07634_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16958_ net253 _01284_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15909_ CPU.registerFile\[18\]\[14\] _03068_ _03069_ CPU.registerFile\[19\]\[14\]
+ _03074_ VGND VGND VPWR VPWR _03394_ sky130_fd_sc_hd__o221a_1
X_16889_ _04169_ VGND VGND VPWR VPWR _04170_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09430_ mapped_spi_ram.rcv_data\[21\] _04688_ _04709_ mapped_spi_flash.rcv_data\[21\]
+ VGND VGND VPWR VPWR _05132_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09361_ net1677 _05066_ _04983_ VGND VGND VPWR VPWR _05067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09292_ _04827_ _04828_ _04905_ VGND VGND VPWR VPWR _05001_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_12 _02856_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 _02940_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_34 _03139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_45 _04730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_56 _04981_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_67 _05093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_78 _05187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_89 _05305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__08468_ clknet_0__08468_ VGND VGND VPWR VPWR clknet_1_1__leaf__08468_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__03970_ clknet_0__03970_ VGND VGND VPWR VPWR clknet_1_0__leaf__03970_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_145_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap14 _04985_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09628_ _04282_ _04806_ VGND VGND VPWR VPWR _05322_ sky130_fd_sc_hd__nor2_1
X_14696__800 clknet_1_1__leaf__02685_ VGND VGND VPWR VPWR net832 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13989__271 clknet_1_1__leaf__08359_ VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_48_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09559_ _04504_ _04647_ _04649_ _04681_ _04654_ VGND VGND VPWR VPWR _05255_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12570_ _07108_ VGND VGND VPWR VPWR _01274_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11521_ net1332 VGND VGND VPWR VPWR _06483_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11452_ _06442_ VGND VGND VPWR VPWR _01797_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10403_ _05830_ _05831_ VGND VGND VPWR VPWR _05832_ sky130_fd_sc_hd__and2_1
X_14171_ CPU.Bimm\[8\] _04718_ _08413_ VGND VGND VPWR VPWR _08423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11383_ _05507_ net1795 _06397_ VGND VGND VPWR VPWR _06406_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13122_ _07291_ _07558_ VGND VGND VPWR VPWR _07559_ sky130_fd_sc_hd__or2_1
X_10334_ _05776_ VGND VGND VPWR VPWR _05788_ sky130_fd_sc_hd__buf_4
XFILLER_0_103_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13053_ _04938_ VGND VGND VPWR VPWR _07492_ sky130_fd_sc_hd__buf_6
X_17930_ net1119 _02214_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_76_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10265_ _05739_ VGND VGND VPWR VPWR _05751_ sky130_fd_sc_hd__clkbuf_4
X_12004_ _05209_ net2065 _06769_ VGND VGND VPWR VPWR _06771_ sky130_fd_sc_hd__mux2_1
X_17861_ net1050 _02145_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_10196_ net2382 _05706_ _05692_ VGND VGND VPWR VPWR _05707_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_880 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16812_ per_uart.uart0.tx_count16\[1\] per_uart.uart0.tx_count16\[0\] VGND VGND VPWR
+ VPWR _04117_ sky130_fd_sc_hd__nand2_1
X_17792_ net981 _02076_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16743_ _04027_ _04039_ _05125_ VGND VGND VPWR VPWR _04062_ sky130_fd_sc_hd__a21o_1
X_12906_ _07238_ VGND VGND VPWR VPWR _07348_ sky130_fd_sc_hd__buf_4
X_16674_ _03998_ _04003_ _06030_ VGND VGND VPWR VPWR _02583_ sky130_fd_sc_hd__a21oi_1
X_13886_ CPU.registerFile\[21\]\[30\] _07502_ _07503_ CPU.registerFile\[17\]\[30\]
+ _07300_ VGND VGND VPWR VPWR _08299_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_17_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15625_ _05070_ VGND VGND VPWR VPWR _03117_ sky130_fd_sc_hd__buf_2
XFILLER_0_9_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12837_ _07273_ _07275_ _07279_ VGND VGND VPWR VPWR _07280_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18344_ clknet_leaf_6_clk _02624_ VGND VGND VPWR VPWR per_uart.rx_error sky130_fd_sc_hd__dfxtp_1
X_15556_ _05405_ VGND VGND VPWR VPWR _03050_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_84_675 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14507_ clknet_1_1__leaf__02664_ VGND VGND VPWR VPWR _02667_ sky130_fd_sc_hd__buf_1
X_11719_ net1444 _06576_ VGND VGND VPWR VPWR _06614_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18275_ net108 _02555_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_15487_ CPU.registerFile\[1\]\[3\] _02814_ _02982_ _02943_ VGND VGND VPWR VPWR _02983_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12699_ per_uart.uart0.enable16_counter\[2\] _07180_ VGND VGND VPWR VPWR _07181_
+ sky130_fd_sc_hd__or2_1
X_17226_ net416 _01514_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__03964_ _03964_ VGND VGND VPWR VPWR clknet_0__03964_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_126_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17157_ net381 _01445_ VGND VGND VPWR VPWR CPU.aluReg\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold805 CPU.registerFile\[15\]\[22\] VGND VGND VPWR VPWR net2046 sky130_fd_sc_hd__dlygate4sd3_1
Xhold816 CPU.registerFile\[31\]\[6\] VGND VGND VPWR VPWR net2057 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16108_ _02924_ _03584_ _03585_ _03586_ _02782_ VGND VGND VPWR VPWR _03587_ sky130_fd_sc_hd__a221o_1
Xhold827 CPU.registerFile\[15\]\[28\] VGND VGND VPWR VPWR net2068 sky130_fd_sc_hd__dlygate4sd3_1
Xhold838 CPU.registerFile\[29\]\[23\] VGND VGND VPWR VPWR net2079 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__02746_ clknet_0__02746_ VGND VGND VPWR VPWR clknet_1_1__leaf__02746_
+ sky130_fd_sc_hd__clkbuf_16
X_17088_ net346 _01410_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[18\] sky130_fd_sc_hd__dfxtp_1
Xhold849 CPU.registerFile\[22\]\[14\] VGND VGND VPWR VPWR net2090 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16039_ CPU.registerFile\[1\]\[18\] _02939_ _03519_ _02894_ VGND VGND VPWR VPWR _03520_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08930_ _04487_ _04624_ VGND VGND VPWR VPWR _04650_ sky130_fd_sc_hd__and2_1
Xclkbuf_1_1__f__02677_ clknet_0__02677_ VGND VGND VPWR VPWR clknet_1_1__leaf__02677_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08861_ _04578_ _04496_ _04458_ _04580_ VGND VGND VPWR VPWR _04581_ sky130_fd_sc_hd__a31o_1
X_08792_ CPU.aluIn1\[9\] CPU.Bimm\[9\] VGND VGND VPWR VPWR _04512_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_127_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14645__754 clknet_1_1__leaf__02680_ VGND VGND VPWR VPWR net786 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_127_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_150_Left_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09413_ _04329_ _04682_ VGND VGND VPWR VPWR _05116_ sky130_fd_sc_hd__nor2_1
X_09344_ _05049_ VGND VGND VPWR VPWR _05050_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_75_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09275_ _04984_ VGND VGND VPWR VPWR _02571_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_43_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14691__796 clknet_1_1__leaf__02684_ VGND VGND VPWR VPWR net828 sky130_fd_sc_hd__inv_2
XFILLER_0_15_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14390__524 clknet_1_1__leaf__02655_ VGND VGND VPWR VPWR net556 sky130_fd_sc_hd__inv_2
XFILLER_0_120_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14728__829 clknet_1_1__leaf__02688_ VGND VGND VPWR VPWR net861 sky130_fd_sc_hd__inv_2
X_10050_ _05620_ VGND VGND VPWR VPWR _02392_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16637__82 clknet_1_1__leaf__03988_ VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__inv_2
XFILLER_0_98_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13740_ _07392_ _08150_ _08157_ VGND VGND VPWR VPWR _08158_ sky130_fd_sc_hd__and3_1
X_10952_ _06176_ VGND VGND VPWR VPWR _02031_ sky130_fd_sc_hd__clkbuf_1
X_16652__96 clknet_1_1__leaf__03989_ VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__inv_2
XFILLER_0_98_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13671_ _07392_ _08088_ _08090_ _07305_ VGND VGND VPWR VPWR _08091_ sky130_fd_sc_hd__a31o_1
X_10883_ _06139_ VGND VGND VPWR VPWR _02063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15410_ CPU.registerFile\[14\]\[2\] CPU.registerFile\[10\]\[2\] _02906_ VGND VGND
+ VPWR VPWR _02907_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__02697_ clknet_0__02697_ VGND VGND VPWR VPWR clknet_1_0__leaf__02697_
+ sky130_fd_sc_hd__clkbuf_16
X_12622_ _07123_ CPU.state\[0\] _07134_ _07135_ VGND VGND VPWR VPWR _00013_ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16390_ _03853_ _03860_ _02844_ VGND VGND VPWR VPWR _03861_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_158_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__07224_ clknet_0__07224_ VGND VGND VPWR VPWR clknet_1_0__leaf__07224_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15341_ CPU.registerFile\[16\]\[0\] _02833_ _02836_ CPU.registerFile\[17\]\[0\] _02764_
+ VGND VGND VPWR VPWR _02840_ sky130_fd_sc_hd__o221a_1
X_12553_ _07099_ VGND VGND VPWR VPWR _01282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18060_ net1233 _02340_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_11504_ _04783_ _06468_ _06470_ VGND VGND VPWR VPWR _06471_ sky130_fd_sc_hd__a21boi_2
X_15272_ _02770_ VGND VGND VPWR VPWR _02771_ sky130_fd_sc_hd__clkbuf_4
X_12484_ net1975 _05696_ _07060_ VGND VGND VPWR VPWR _07063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17011_ net269 _01333_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_78_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11435_ _05487_ net2402 _06433_ VGND VGND VPWR VPWR _06434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__02700_ _02700_ VGND VGND VPWR VPWR clknet_0__02700_ sky130_fd_sc_hd__clkbuf_16
X_14154_ CPU.Iimm\[0\] _07653_ _08413_ VGND VGND VPWR VPWR _08414_ sky130_fd_sc_hd__mux2_1
X_11366_ _06396_ VGND VGND VPWR VPWR _06397_ sky130_fd_sc_hd__buf_4
XFILLER_0_21_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13105_ CPU.registerFile\[2\]\[6\] CPU.registerFile\[3\]\[6\] _07260_ VGND VGND VPWR
+ VPWR _07542_ sky130_fd_sc_hd__mux2_1
X_10317_ _05779_ VGND VGND VPWR VPWR _02269_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_91_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11297_ _06359_ VGND VGND VPWR VPWR _06360_ sky130_fd_sc_hd__buf_4
X_13036_ _07296_ VGND VGND VPWR VPWR _07475_ sky130_fd_sc_hd__buf_4
X_10248_ _05742_ VGND VGND VPWR VPWR _02316_ sky130_fd_sc_hd__clkbuf_1
X_17913_ net1102 net1317 VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14367__504 clknet_1_0__leaf__02652_ VGND VGND VPWR VPWR net536 sky130_fd_sc_hd__inv_2
X_17844_ net1033 _02128_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_10179_ _05695_ VGND VGND VPWR VPWR _02338_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_109_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17775_ net964 _02059_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_16726_ _08457_ _04045_ _04046_ _04047_ VGND VGND VPWR VPWR _04048_ sky130_fd_sc_hd__a31o_1
X_13938_ CPU.registerFile\[30\]\[31\] CPU.registerFile\[26\]\[31\] _04937_ VGND VGND
+ VPWR VPWR _08350_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_122_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13869_ _07818_ _08281_ _08282_ VGND VGND VPWR VPWR _08283_ sky130_fd_sc_hd__o21a_1
XFILLER_0_158_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15608_ CPU.registerFile\[5\]\[6\] CPU.registerFile\[4\]\[6\] _02805_ VGND VGND VPWR
+ VPWR _03101_ sky130_fd_sc_hd__mux2_1
X_16588_ clknet_1_1__leaf__07219_ VGND VGND VPWR VPWR _03970_ sky130_fd_sc_hd__buf_1
XFILLER_0_45_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18327_ clknet_leaf_6_clk _02607_ VGND VGND VPWR VPWR per_uart.uart0.tx_count16\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15539_ _03030_ _03031_ _03033_ _02901_ VGND VGND VPWR VPWR _03034_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09060_ _04769_ _04770_ _04772_ _04773_ VGND VGND VPWR VPWR _04774_ sky130_fd_sc_hd__o31a_1
XFILLER_0_60_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18258_ net99 _02538_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17209_ net399 _01497_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_18189_ net220 _02469_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[23\] sky130_fd_sc_hd__dfxtp_1
Xhold602 per_uart.uart0.txd_reg\[5\] VGND VGND VPWR VPWR net1843 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold613 CPU.registerFile\[27\]\[18\] VGND VGND VPWR VPWR net1854 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold624 CPU.registerFile\[3\]\[22\] VGND VGND VPWR VPWR net1865 sky130_fd_sc_hd__dlygate4sd3_1
Xhold635 CPU.registerFile\[23\]\[0\] VGND VGND VPWR VPWR net1876 sky130_fd_sc_hd__dlygate4sd3_1
Xhold646 CPU.registerFile\[21\]\[17\] VGND VGND VPWR VPWR net1887 sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 CPU.registerFile\[18\]\[15\] VGND VGND VPWR VPWR net1898 sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 CPU.registerFile\[1\]\[9\] VGND VGND VPWR VPWR net1909 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09962_ _05573_ VGND VGND VPWR VPWR _02465_ sky130_fd_sc_hd__clkbuf_1
Xhold679 CPU.registerFile\[18\]\[21\] VGND VGND VPWR VPWR net1920 sky130_fd_sc_hd__dlygate4sd3_1
X_15240__149 clknet_1_0__leaf__02754_ VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__inv_2
X_08913_ _04520_ _04632_ _04590_ VGND VGND VPWR VPWR _04633_ sky130_fd_sc_hd__o21a_1
X_09893_ _05169_ VGND VGND VPWR VPWR _05530_ sky130_fd_sc_hd__clkbuf_8
Xhold1302 mapped_spi_flash.snd_bitcount\[2\] VGND VGND VPWR VPWR net2543 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08844_ _04563_ _04562_ VGND VGND VPWR VPWR _04564_ sky130_fd_sc_hd__or2_4
X_08775_ _04494_ VGND VGND VPWR VPWR _04495_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09327_ _04252_ _04336_ VGND VGND VPWR VPWR _05034_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09258_ _04245_ _04214_ _04965_ _04967_ VGND VGND VPWR VPWR _04968_ sky130_fd_sc_hd__a211o_1
XFILLER_0_63_678 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_153_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09189_ _04843_ _04899_ _04900_ VGND VGND VPWR VPWR _04901_ sky130_fd_sc_hd__o21ai_1
X_11220_ _05549_ net2192 _06310_ VGND VGND VPWR VPWR _06319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14972__1049 clknet_1_0__leaf__02712_ VGND VGND VPWR VPWR net1081 sky130_fd_sc_hd__inv_2
X_11151_ _06282_ VGND VGND VPWR VPWR _01938_ sky130_fd_sc_hd__clkbuf_1
X_14316__458 clknet_1_1__leaf__08464_ VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_56_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10102_ _05648_ VGND VGND VPWR VPWR _02368_ sky130_fd_sc_hd__clkbuf_1
X_11082_ _06245_ VGND VGND VPWR VPWR _01970_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_8_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10033_ _05611_ VGND VGND VPWR VPWR _02400_ sky130_fd_sc_hd__clkbuf_1
X_15890_ CPU.registerFile\[30\]\[14\] CPU.registerFile\[26\]\[14\] _03247_ VGND VGND
+ VPWR VPWR _03375_ sky130_fd_sc_hd__mux2_1
X_17560_ net749 _01848_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_11984_ _06760_ VGND VGND VPWR VPWR _01580_ sky130_fd_sc_hd__clkbuf_1
X_16511_ clknet_1_0__leaf__02749_ VGND VGND VPWR VPWR _03963_ sky130_fd_sc_hd__buf_1
XFILLER_0_98_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13723_ net1480 _08018_ _08141_ _08017_ VGND VGND VPWR VPWR _01319_ sky130_fd_sc_hd__o211a_1
X_10935_ net1579 _05717_ _06165_ VGND VGND VPWR VPWR _06168_ sky130_fd_sc_hd__mux2_1
X_17491_ net680 _01779_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[5\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_104_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__02749_ clknet_0__02749_ VGND VGND VPWR VPWR clknet_1_0__leaf__02749_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_27_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16442_ _03904_ _03910_ _02879_ VGND VGND VPWR VPWR _03911_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_27_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13654_ _07245_ _08074_ VGND VGND VPWR VPWR _08075_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10866_ net2339 _05717_ _06128_ VGND VGND VPWR VPWR _06131_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12605_ _05820_ _05819_ VGND VGND VPWR VPWR _07125_ sky130_fd_sc_hd__nor2_1
X_16373_ CPU.registerFile\[29\]\[28\] _02918_ VGND VGND VPWR VPWR _03844_ sky130_fd_sc_hd__or2_1
X_13585_ _07291_ _08007_ VGND VGND VPWR VPWR _08008_ sky130_fd_sc_hd__or2_1
X_10797_ _06094_ VGND VGND VPWR VPWR _02104_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18112_ net175 _02392_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[10\] sky130_fd_sc_hd__dfxtp_1
X_15324_ CPU.registerFile\[2\]\[0\] _02821_ _02822_ CPU.registerFile\[3\]\[0\] _05070_
+ VGND VGND VPWR VPWR _02823_ sky130_fd_sc_hd__a221o_1
XFILLER_0_54_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12536_ _07090_ VGND VGND VPWR VPWR _01290_ sky130_fd_sc_hd__clkbuf_1
X_14674__780 clknet_1_1__leaf__02683_ VGND VGND VPWR VPWR net812 sky130_fd_sc_hd__inv_2
XFILLER_0_30_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18043_ net1216 _02323_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12467_ net1874 _05679_ _07049_ VGND VGND VPWR VPWR _07054_ sky130_fd_sc_hd__mux2_1
XFILLER_0_112_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_144_Right_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11418_ _06424_ VGND VGND VPWR VPWR _01813_ sky130_fd_sc_hd__clkbuf_1
X_15186_ clknet_1_1__leaf__02749_ VGND VGND VPWR VPWR _02750_ sky130_fd_sc_hd__buf_1
X_12398_ _07017_ VGND VGND VPWR VPWR _01388_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14137_ _08400_ VGND VGND VPWR VPWR _08401_ sky130_fd_sc_hd__buf_4
X_11349_ _06387_ VGND VGND VPWR VPWR _01845_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14072__346 clknet_1_0__leaf__08367_ VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__inv_2
X_13019_ CPU.registerFile\[18\]\[4\] CPU.registerFile\[22\]\[4\] _07457_ VGND VGND
+ VPWR VPWR _07458_ sky130_fd_sc_hd__mux2_1
X_17827_ net1016 _02111_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08560_ CPU.aluIn1\[5\] _04279_ VGND VGND VPWR VPWR _04280_ sky130_fd_sc_hd__nand2_1
X_17758_ net947 _02042_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08491_ _04210_ VGND VGND VPWR VPWR _04211_ sky130_fd_sc_hd__clkbuf_4
X_16709_ _04032_ CPU.PC\[9\] VGND VGND VPWR VPWR _04033_ sky130_fd_sc_hd__and2_1
X_17689_ net878 _01977_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_16631__77 clknet_1_1__leaf__03971_ VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__inv_2
XFILLER_0_9_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14757__855 clknet_1_0__leaf__02691_ VGND VGND VPWR VPWR net887 sky130_fd_sc_hd__inv_2
XFILLER_0_147_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16517__185 clknet_1_1__leaf__03963_ VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_40_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09112_ CPU.PC\[21\] _04822_ VGND VGND VPWR VPWR _04824_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09043_ mapped_spi_ram.rcv_data\[2\] _04689_ _04691_ mapped_spi_flash.rcv_data\[2\]
+ VGND VGND VPWR VPWR _04758_ sky130_fd_sc_hd__a22o_2
XFILLER_0_143_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_135_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold410 CPU.registerFile\[14\]\[26\] VGND VGND VPWR VPWR net1651 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_111_Right_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold421 CPU.registerFile\[28\]\[30\] VGND VGND VPWR VPWR net1662 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold432 CPU.registerFile\[5\]\[0\] VGND VGND VPWR VPWR net1673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 per_uart.uart0.rx_bitcount\[3\] VGND VGND VPWR VPWR net1684 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold454 CPU.registerFile\[18\]\[20\] VGND VGND VPWR VPWR net1695 sky130_fd_sc_hd__dlygate4sd3_1
Xhold465 CPU.registerFile\[16\]\[31\] VGND VGND VPWR VPWR net1706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 CPU.registerFile\[16\]\[21\] VGND VGND VPWR VPWR net1717 sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 CPU.registerFile\[29\]\[24\] VGND VGND VPWR VPWR net1728 sky130_fd_sc_hd__dlygate4sd3_1
Xhold498 CPU.registerFile\[7\]\[31\] VGND VGND VPWR VPWR net1739 sky130_fd_sc_hd__dlygate4sd3_1
X_09945_ _05564_ VGND VGND VPWR VPWR _02473_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ _05518_ net2440 _05512_ VGND VGND VPWR VPWR _05519_ sky130_fd_sc_hd__mux2_1
Xhold1110 CPU.registerFile\[19\]\[22\] VGND VGND VPWR VPWR net2351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1121 CPU.registerFile\[21\]\[5\] VGND VGND VPWR VPWR net2362 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1132 CPU.registerFile\[27\]\[7\] VGND VGND VPWR VPWR net2373 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ _04543_ _04512_ _04544_ _04546_ VGND VGND VPWR VPWR _04547_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_51_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1143 CPU.rs2\[8\] VGND VGND VPWR VPWR net2384 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1154 CPU.registerFile\[21\]\[6\] VGND VGND VPWR VPWR net2395 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1165 CPU.registerFile\[15\]\[16\] VGND VGND VPWR VPWR net2406 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1176 CPU.registerFile\[28\]\[19\] VGND VGND VPWR VPWR net2417 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1187 CPU.rs2\[10\] VGND VGND VPWR VPWR net2428 sky130_fd_sc_hd__dlygate4sd3_1
X_08758_ _04378_ _04477_ _04367_ VGND VGND VPWR VPWR _04478_ sky130_fd_sc_hd__o21ba_1
XANTENNA_305 _07412_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1198 mapped_spi_ram.snd_bitcount\[5\] VGND VGND VPWR VPWR net2439 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_316 _07914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_327 _07953_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_338 _02895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08689_ _04297_ _04299_ VGND VGND VPWR VPWR _04409_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_349 _05380_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10720_ _06053_ VGND VGND VPWR VPWR _02140_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_24_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10651_ mapped_spi_flash.div_counter\[0\] net1314 VGND VGND VPWR VPWR _06011_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13370_ _07584_ _07784_ _07799_ _07309_ VGND VGND VPWR VPWR _07800_ sky130_fd_sc_hd__a211o_1
X_10582_ net1453 _05968_ _05972_ _05936_ VGND VGND VPWR VPWR _02196_ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12321_ _05775_ _06032_ VGND VGND VPWR VPWR _06976_ sky130_fd_sc_hd__nand2_2
XFILLER_0_121_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12252_ _06861_ VGND VGND VPWR VPWR _06924_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11203_ _06287_ VGND VGND VPWR VPWR _06310_ sky130_fd_sc_hd__buf_4
X_12183_ _04483_ _05134_ VGND VGND VPWR VPWR _06870_ sky130_fd_sc_hd__nor2_1
X_15223__133 clknet_1_0__leaf__02753_ VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_71_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11134_ _06273_ VGND VGND VPWR VPWR _01946_ sky130_fd_sc_hd__clkbuf_1
X_16991_ clknet_leaf_21_clk _01317_ VGND VGND VPWR VPWR CPU.rs2\[22\] sky130_fd_sc_hd__dfxtp_1
X_11065_ _06236_ VGND VGND VPWR VPWR _01978_ sky130_fd_sc_hd__clkbuf_1
X_15942_ CPU.registerFile\[19\]\[15\] CPU.registerFile\[17\]\[15\] _02874_ VGND VGND
+ VPWR VPWR _03426_ sky130_fd_sc_hd__mux2_1
X_10016_ _05602_ VGND VGND VPWR VPWR _02408_ sky130_fd_sc_hd__clkbuf_1
X_15873_ _03065_ _03357_ _03358_ VGND VGND VPWR VPWR _03359_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17612_ net801 _01900_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_17543_ net732 _01831_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11967_ _06751_ VGND VGND VPWR VPWR _01588_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14479__605 clknet_1_0__leaf__02663_ VGND VGND VPWR VPWR net637 sky130_fd_sc_hd__inv_2
X_13706_ _08121_ _08124_ _07514_ VGND VGND VPWR VPWR _08125_ sky130_fd_sc_hd__a21oi_4
X_10918_ net1573 _05700_ _06154_ VGND VGND VPWR VPWR _06159_ sky130_fd_sc_hd__mux2_1
X_17474_ net663 _01762_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[29\] sky130_fd_sc_hd__dfxtp_1
X_11898_ net2424 _05677_ _06711_ VGND VGND VPWR VPWR _06715_ sky130_fd_sc_hd__mux2_1
X_16425_ _03890_ _03894_ _02810_ VGND VGND VPWR VPWR _03895_ sky130_fd_sc_hd__a21o_1
XFILLER_0_129_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13637_ CPU.registerFile\[21\]\[22\] _07361_ _07283_ CPU.registerFile\[17\]\[22\]
+ _07554_ VGND VGND VPWR VPWR _08058_ sky130_fd_sc_hd__o221a_1
X_10849_ net1970 _05700_ _06117_ VGND VGND VPWR VPWR _06122_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_128_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16356_ _02903_ _03818_ _03827_ _03252_ VGND VGND VPWR VPWR _03828_ sky130_fd_sc_hd__o211a_1
X_13568_ CPU.registerFile\[5\]\[20\] _07804_ _07990_ _07368_ VGND VGND VPWR VPWR _07991_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15307_ _02805_ VGND VGND VPWR VPWR _02806_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12519_ net1929 _05731_ _07071_ VGND VGND VPWR VPWR _07081_ sky130_fd_sc_hd__mux2_1
X_16287_ _02858_ _03757_ _03760_ _02809_ VGND VGND VPWR VPWR _03761_ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13499_ _07364_ _07923_ VGND VGND VPWR VPWR _07924_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_117_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18026_ net1199 _02306_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15198__110 clknet_1_1__leaf__02751_ VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_130_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09730_ _04672_ _05416_ _05419_ _04679_ VGND VGND VPWR VPWR _05420_ sky130_fd_sc_hd__o211a_1
XFILLER_0_66_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09661_ _05351_ _05353_ _04670_ VGND VGND VPWR VPWR _05354_ sky130_fd_sc_hd__mux2_1
X_08612_ _04331_ VGND VGND VPWR VPWR _04332_ sky130_fd_sc_hd__inv_2
X_09592_ _05275_ _05276_ _05285_ _05286_ VGND VGND VPWR VPWR _05287_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_19_Left_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08543_ CPU.rs2\[10\] CPU.Bimm\[10\] net1295 VGND VGND VPWR VPWR _04263_ sky130_fd_sc_hd__mux2_1
X_14971__1048 clknet_1_0__leaf__02712_ VGND VGND VPWR VPWR net1080 sky130_fd_sc_hd__inv_2
XFILLER_0_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14345__484 clknet_1_1__leaf__08467_ VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__inv_2
XFILLER_0_148_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08474_ mapped_spi_ram.div_counter\[0\] mapped_spi_ram.div_counter\[1\] net23 _04193_
+ VGND VGND VPWR VPWR _04195_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_9_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13983__266 clknet_1_0__leaf__08358_ VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__inv_2
XFILLER_0_135_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_150_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_28_Left_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09026_ _04230_ _04698_ _04218_ CPU.aluReg\[27\] _04741_ VGND VGND VPWR VPWR _04742_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold240 mapped_spi_ram.rcv_data\[6\] VGND VGND VPWR VPWR net1481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 CPU.cycles\[1\] VGND VGND VPWR VPWR net1492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 mapped_spi_ram.rcv_data\[18\] VGND VGND VPWR VPWR net1503 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 CPU.cycles\[13\] VGND VGND VPWR VPWR net1514 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14055__330 clknet_1_0__leaf__08366_ VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__inv_2
XFILLER_0_130_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold284 CPU.cycles\[7\] VGND VGND VPWR VPWR net1525 sky130_fd_sc_hd__dlygate4sd3_1
X_14510__632 clknet_1_1__leaf__02667_ VGND VGND VPWR VPWR net664 sky130_fd_sc_hd__inv_2
Xhold295 per_uart.uart_ctrl\[2\] VGND VGND VPWR VPWR net1536 sky130_fd_sc_hd__dlygate4sd3_1
X_09928_ _05553_ net2025 _05490_ VGND VGND VPWR VPWR _05554_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_148_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_148_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09859_ _04932_ VGND VGND VPWR VPWR _05507_ sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_37_Left_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14428__559 clknet_1_1__leaf__02658_ VGND VGND VPWR VPWR net591 sky130_fd_sc_hd__inv_2
X_12870_ CPU.registerFile\[2\]\[1\] CPU.registerFile\[3\]\[1\] _07311_ VGND VGND VPWR
+ VPWR _07312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_102 _05381_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11821_ _06673_ VGND VGND VPWR VPWR _01656_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_113 _05426_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_124 _05530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_135 _05694_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_146 _07260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_157 _07291_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14540_ clknet_1_0__leaf__02664_ VGND VGND VPWR VPWR _02670_ sky130_fd_sc_hd__buf_1
XANTENNA_168 _07330_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11752_ _06637_ VGND VGND VPWR VPWR _01689_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_179 _07507_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10703_ _06044_ VGND VGND VPWR VPWR _02148_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11683_ net1503 _06590_ _06593_ _06594_ VGND VGND VPWR VPWR _01714_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_81_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16210_ _02796_ _03685_ VGND VGND VPWR VPWR _03686_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_81_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13422_ CPU.registerFile\[15\]\[15\] _07276_ _07277_ CPU.registerFile\[11\]\[15\]
+ _07820_ VGND VGND VPWR VPWR _07850_ sky130_fd_sc_hd__o221a_1
XFILLER_0_64_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17190_ clknet_leaf_25_clk _01478_ VGND VGND VPWR VPWR CPU.Iimm\[0\] sky130_fd_sc_hd__dfxtp_2
X_10634_ net1506 _05996_ _06001_ _05993_ VGND VGND VPWR VPWR _02173_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16141_ CPU.registerFile\[2\]\[21\] _03143_ _02980_ CPU.registerFile\[3\]\[21\] _03144_
+ VGND VGND VPWR VPWR _03619_ sky130_fd_sc_hd__a221o_1
X_13353_ _07780_ _07782_ _07320_ VGND VGND VPWR VPWR _07783_ sky130_fd_sc_hd__mux2_1
X_10565_ net1507 net2544 VGND VGND VPWR VPWR _05959_ sky130_fd_sc_hd__nor2_1
X_12304_ _06963_ VGND VGND VPWR VPWR _01428_ sky130_fd_sc_hd__clkbuf_1
X_16072_ CPU.registerFile\[13\]\[19\] _02775_ VGND VGND VPWR VPWR _03552_ sky130_fd_sc_hd__or2_1
X_13284_ CPU.registerFile\[21\]\[11\] _07362_ _07363_ CPU.registerFile\[17\]\[11\]
+ _07715_ VGND VGND VPWR VPWR _07716_ sky130_fd_sc_hd__o221a_2
X_10496_ _05903_ _04544_ _04543_ VGND VGND VPWR VPWR _05904_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_121_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12235_ CPU.aluIn1\[20\] _06910_ _06894_ VGND VGND VPWR VPWR _06911_ sky130_fd_sc_hd__mux2_1
X_14786__881 clknet_1_0__leaf__02694_ VGND VGND VPWR VPWR net913 sky130_fd_sc_hd__inv_2
X_12166_ CPU.aluShamt\[4\] _06854_ VGND VGND VPWR VPWR _06858_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_112_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11117_ CPU.registerFile\[8\]\[20\] _05694_ _06263_ VGND VGND VPWR VPWR _06265_ sky130_fd_sc_hd__mux2_1
X_16974_ clknet_leaf_22_clk _01300_ VGND VGND VPWR VPWR CPU.mem_wdata\[5\] sky130_fd_sc_hd__dfxtp_2
X_12097_ _06820_ VGND VGND VPWR VPWR _01526_ sky130_fd_sc_hd__clkbuf_1
X_15925_ CPU.registerFile\[6\]\[15\] CPU.registerFile\[7\]\[15\] _02870_ VGND VGND
+ VPWR VPWR _03409_ sky130_fd_sc_hd__mux2_1
X_11048_ CPU.registerFile\[7\]\[20\] _05694_ _06226_ VGND VGND VPWR VPWR _06228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15856_ CPU.registerFile\[30\]\[13\] CPU.registerFile\[26\]\[13\] _02787_ VGND VGND
+ VPWR VPWR _03342_ sky130_fd_sc_hd__mux2_1
X_15787_ CPU.registerFile\[28\]\[11\] _02791_ VGND VGND VPWR VPWR _03275_ sky130_fd_sc_hd__or2_1
X_12999_ _04939_ _07436_ _07438_ _04972_ VGND VGND VPWR VPWR _07439_ sky130_fd_sc_hd__a211o_1
XFILLER_0_98_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14225__400 clknet_1_0__leaf__08432_ VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__inv_2
XFILLER_0_87_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17526_ net715 _01814_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_578 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17457_ net646 _01745_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_119_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16408_ CPU.registerFile\[8\]\[29\] CPU.registerFile\[12\]\[29\] _03254_ VGND VGND
+ VPWR VPWR _03878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17388_ net577 _01676_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16339_ CPU.registerFile\[22\]\[27\] _05049_ VGND VGND VPWR VPWR _03811_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_732 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14869__956 clknet_1_1__leaf__02702_ VGND VGND VPWR VPWR net988 sky130_fd_sc_hd__inv_2
XFILLER_0_152_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18009_ net1182 _02289_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09713_ _05403_ VGND VGND VPWR VPWR _02552_ sky130_fd_sc_hd__clkbuf_1
X_09644_ _05336_ VGND VGND VPWR VPWR _05337_ sky130_fd_sc_hd__buf_4
XFILLER_0_93_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09575_ _04651_ _05255_ _05270_ VGND VGND VPWR VPWR _05271_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_143_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08526_ CPU.rs2\[20\] _04200_ _04205_ VGND VGND VPWR VPWR _04246_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_795 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10350_ _05796_ VGND VGND VPWR VPWR _02253_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09009_ _04363_ _04670_ _04725_ VGND VGND VPWR VPWR _04726_ sky130_fd_sc_hd__and3b_1
XFILLER_0_60_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10281_ _05759_ VGND VGND VPWR VPWR _02300_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12020_ _05402_ net1904 _06769_ VGND VGND VPWR VPWR _06779_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_45_Left_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15710_ _08397_ _03194_ _03199_ _02903_ VGND VGND VPWR VPWR _03200_ sky130_fd_sc_hd__o211a_1
X_12922_ _07283_ VGND VGND VPWR VPWR _07363_ sky130_fd_sc_hd__clkbuf_8
X_16690_ _08436_ _08459_ _05293_ VGND VGND VPWR VPWR _04017_ sky130_fd_sc_hd__a21oi_1
X_15641_ _02786_ _03129_ _03132_ _02794_ VGND VGND VPWR VPWR _03133_ sky130_fd_sc_hd__a211o_1
XFILLER_0_87_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12853_ _05338_ VGND VGND VPWR VPWR _07296_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_158_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ _05253_ net2175 _06661_ VGND VGND VPWR VPWR _06665_ sky130_fd_sc_hd__mux2_1
X_18360_ clknet_leaf_5_clk _02638_ VGND VGND VPWR VPWR per_uart.d_in_uart\[0\] sky130_fd_sc_hd__dfxtp_1
X_15572_ _08394_ VGND VGND VPWR VPWR _03066_ sky130_fd_sc_hd__buf_4
XFILLER_0_84_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12784_ CPU.state\[2\] _07120_ VGND VGND VPWR VPWR _07227_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17311_ net500 _01599_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_835 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13966__250 clknet_1_0__leaf__08357_ VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__inv_2
XFILLER_0_113_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18291_ net124 _02571_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_11735_ _06572_ _06569_ net2 VGND VGND VPWR VPWR _00008_ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_54_Left_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17242_ net432 _01530_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11666_ net1322 _06575_ _06584_ _06581_ VGND VGND VPWR VPWR _01721_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_12_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13405_ _07230_ _07817_ _07833_ _07309_ VGND VGND VPWR VPWR _07834_ sky130_fd_sc_hd__a211o_1
X_17173_ clknet_leaf_12_clk _01461_ VGND VGND VPWR VPWR CPU.instr\[3\] sky130_fd_sc_hd__dfxtp_2
X_10617_ mapped_spi_flash.rcv_data\[13\] _05983_ _05991_ _05980_ VGND VGND VPWR VPWR
+ _02180_ sky130_fd_sc_hd__o211a_1
X_14385_ clknet_1_0__leaf__02653_ VGND VGND VPWR VPWR _02655_ sky130_fd_sc_hd__buf_1
XFILLER_0_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11597_ net1359 _06524_ _06536_ _06516_ VGND VGND VPWR VPWR _01742_ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16124_ _02786_ _03599_ _03601_ _03019_ VGND VGND VPWR VPWR _03602_ sky130_fd_sc_hd__a211o_1
XFILLER_0_12_607 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13336_ _07271_ _07755_ _07758_ _07765_ _07766_ VGND VGND VPWR VPWR _07767_ sky130_fd_sc_hd__o311a_1
X_14220__396 clknet_1_1__leaf__08431_ VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_114_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10548_ mapped_spi_flash.snd_bitcount\[5\] _05945_ VGND VGND VPWR VPWR _05946_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16055_ CPU.registerFile\[2\]\[19\] _03227_ _03228_ CPU.registerFile\[3\]\[19\] _03534_
+ VGND VGND VPWR VPWR _03535_ sky130_fd_sc_hd__a221o_1
X_13267_ CPU.registerFile\[15\]\[10\] _07402_ _07500_ CPU.registerFile\[11\]\[10\]
+ _07327_ VGND VGND VPWR VPWR _07700_ sky130_fd_sc_hd__o221a_1
Xclkbuf_1_1__f__02693_ clknet_0__02693_ VGND VGND VPWR VPWR clknet_1_1__leaf__02693_
+ sky130_fd_sc_hd__clkbuf_16
X_14970__1047 clknet_1_0__leaf__02712_ VGND VGND VPWR VPWR net1079 sky130_fd_sc_hd__inv_2
X_10479_ _05852_ _05889_ VGND VGND VPWR VPWR _05890_ sky130_fd_sc_hd__nor2_1
X_15006_ clknet_1_1__leaf__02708_ VGND VGND VPWR VPWR _02716_ sky130_fd_sc_hd__buf_1
X_12218_ CPU.aluIn1\[24\] _06897_ _06894_ VGND VGND VPWR VPWR _06898_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__07220_ clknet_0__07220_ VGND VGND VPWR VPWR clknet_1_1__leaf__07220_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_94_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13198_ CPU.registerFile\[31\]\[8\] _07402_ _07500_ CPU.registerFile\[27\]\[8\] _07483_
+ VGND VGND VPWR VPWR _07633_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_63_Left_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12149_ _06847_ VGND VGND VPWR VPWR _01501_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16957_ net252 _01283_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_15908_ CPU.registerFile\[22\]\[14\] CPU.registerFile\[23\]\[14\] _02828_ VGND VGND
+ VPWR VPWR _03393_ sky130_fd_sc_hd__mux2_1
X_16888_ per_uart.uart0.rx_bitcount\[2\] per_uart.uart0.rx_bitcount\[1\] per_uart.uart0.rx_bitcount\[0\]
+ _04164_ _04165_ VGND VGND VPWR VPWR _04169_ sky130_fd_sc_hd__a41o_1
XFILLER_0_78_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15839_ _03065_ _03324_ _03325_ VGND VGND VPWR VPWR _03326_ sky130_fd_sc_hd__o21a_1
XFILLER_0_149_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09360_ _05065_ VGND VGND VPWR VPWR _05066_ sky130_fd_sc_hd__buf_8
XFILLER_0_75_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_72_Left_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_904 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17509_ net698 _01797_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09291_ _04992_ _04999_ _04773_ VGND VGND VPWR VPWR _05000_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_13 _02861_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_24 _02948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_35 _03176_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_46 _04730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_57 _04981_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_68 _05093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_79 _05187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14457__585 clknet_1_1__leaf__02661_ VGND VGND VPWR VPWR net617 sky130_fd_sc_hd__inv_2
XFILLER_0_30_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14195__373 clknet_1_1__leaf__08429_ VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__inv_2
XFILLER_0_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__08467_ clknet_0__08467_ VGND VGND VPWR VPWR clknet_1_1__leaf__08467_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_112_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_81_Left_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_145_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap15 _04620_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_4
X_09627_ _04800_ _05318_ _05320_ _04768_ VGND VGND VPWR VPWR _05321_ sky130_fd_sc_hd__o211a_1
X_14622__733 clknet_1_1__leaf__02678_ VGND VGND VPWR VPWR net765 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_39_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09558_ _05254_ VGND VGND VPWR VPWR _02558_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08509_ CPU.rs2\[27\] _04201_ _04206_ VGND VGND VPWR VPWR _04229_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09489_ _04667_ VGND VGND VPWR VPWR _05189_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_61_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11520_ _04192_ VGND VGND VPWR VPWR _06482_ sky130_fd_sc_hd__buf_4
XFILLER_0_93_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11451_ _05507_ net2276 _06433_ VGND VGND VPWR VPWR _06442_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10402_ mapped_spi_flash.cmd_addr\[29\] _05825_ _05827_ mapped_spi_flash.cmd_addr\[30\]
+ VGND VGND VPWR VPWR _05831_ sky130_fd_sc_hd__a22o_1
X_14170_ _08422_ VGND VGND VPWR VPWR _01485_ sky130_fd_sc_hd__clkbuf_1
X_11382_ _06405_ VGND VGND VPWR VPWR _01830_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13121_ CPU.registerFile\[28\]\[6\] CPU.registerFile\[24\]\[6\] _07292_ VGND VGND
+ VPWR VPWR _07558_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10333_ _05787_ VGND VGND VPWR VPWR _02261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13052_ _07412_ _07487_ _07490_ VGND VGND VPWR VPWR _07491_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_76_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10264_ _05750_ VGND VGND VPWR VPWR _02308_ sky130_fd_sc_hd__clkbuf_1
X_12003_ _06770_ VGND VGND VPWR VPWR _01571_ sky130_fd_sc_hd__clkbuf_1
X_10195_ _05129_ VGND VGND VPWR VPWR _05706_ sky130_fd_sc_hd__clkbuf_4
X_17860_ net1049 _02144_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16811_ net1529 _08355_ _04116_ _03632_ VGND VGND VPWR VPWR _02607_ sky130_fd_sc_hd__o211a_1
X_17791_ net980 _02075_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_916 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13954_ clknet_1_1__leaf__07223_ VGND VGND VPWR VPWR _08356_ sky130_fd_sc_hd__buf_1
X_16742_ _04032_ net1569 VGND VGND VPWR VPWR _04061_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12905_ _07235_ VGND VGND VPWR VPWR _07347_ sky130_fd_sc_hd__buf_4
X_14898__982 clknet_1_1__leaf__02705_ VGND VGND VPWR VPWR net1014 sky130_fd_sc_hd__inv_2
X_16673_ _08457_ _03999_ _04000_ _04002_ VGND VGND VPWR VPWR _04003_ sky130_fd_sc_hd__a31o_1
X_13885_ CPU.registerFile\[23\]\[30\] _07325_ _07500_ CPU.registerFile\[19\]\[30\]
+ _07327_ VGND VGND VPWR VPWR _08298_ sky130_fd_sc_hd__o221a_1
XFILLER_0_69_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14597__710 clknet_1_1__leaf__02676_ VGND VGND VPWR VPWR net742 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15624_ CPU.registerFile\[14\]\[7\] CPU.registerFile\[10\]\[7\] _03082_ VGND VGND
+ VPWR VPWR _03116_ sky130_fd_sc_hd__mux2_1
X_12836_ CPU.registerFile\[15\]\[0\] _07276_ _07277_ CPU.registerFile\[11\]\[0\] _07278_
+ VGND VGND VPWR VPWR _07279_ sky130_fd_sc_hd__o221a_1
XFILLER_0_69_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15555_ _02786_ _03046_ _03048_ _02794_ VGND VGND VPWR VPWR _03049_ sky130_fd_sc_hd__a211o_1
X_18343_ clknet_leaf_5_clk _02623_ VGND VGND VPWR VPWR per_uart.rx_data\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11718_ net1444 _06603_ _06613_ _06607_ VGND VGND VPWR VPWR _01698_ sky130_fd_sc_hd__o211a_1
X_18274_ net107 _02554_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15486_ CPU.registerFile\[5\]\[3\] CPU.registerFile\[4\]\[3\] _02805_ VGND VGND VPWR
+ VPWR _02982_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12698_ net1363 per_uart.uart0.enable16_counter\[0\] VGND VGND VPWR VPWR _07180_
+ sky130_fd_sc_hd__or2_1
Xclkbuf_0__03963_ _03963_ VGND VGND VPWR VPWR clknet_0__03963_ sky130_fd_sc_hd__clkbuf_16
X_17225_ net415 _01513_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_11649_ _06569_ _06572_ VGND VGND VPWR VPWR _06573_ sky130_fd_sc_hd__or2b_1
XFILLER_0_52_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17156_ net380 _01444_ VGND VGND VPWR VPWR CPU.aluReg\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold806 CPU.registerFile\[8\]\[29\] VGND VGND VPWR VPWR net2047 sky130_fd_sc_hd__dlygate4sd3_1
X_16107_ CPU.registerFile\[13\]\[20\] _02775_ VGND VGND VPWR VPWR _03586_ sky130_fd_sc_hd__or2_1
Xhold817 CPU.registerFile\[27\]\[28\] VGND VGND VPWR VPWR net2058 sky130_fd_sc_hd__dlygate4sd3_1
X_13319_ _04939_ _07747_ _07749_ _04972_ VGND VGND VPWR VPWR _07750_ sky130_fd_sc_hd__a211o_1
XFILLER_0_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold828 per_uart.uart0.rxd_reg\[2\] VGND VGND VPWR VPWR net2069 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold839 CPU.registerFile\[13\]\[19\] VGND VGND VPWR VPWR net2080 sky130_fd_sc_hd__dlygate4sd3_1
X_17087_ net345 _01409_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[17\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__02745_ clknet_0__02745_ VGND VGND VPWR VPWR clknet_1_1__leaf__02745_
+ sky130_fd_sc_hd__clkbuf_16
X_16038_ CPU.registerFile\[5\]\[18\] CPU.registerFile\[4\]\[18\] _03146_ VGND VGND
+ VPWR VPWR _03519_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__02676_ clknet_0__02676_ VGND VGND VPWR VPWR clknet_1_1__leaf__02676_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08860_ _04496_ _04579_ CPU.aluIn1\[22\] CPU.aluIn1\[21\] VGND VGND VPWR VPWR _04580_
+ sky130_fd_sc_hd__and4b_1
X_08791_ CPU.aluIn1\[10\] CPU.Bimm\[10\] VGND VGND VPWR VPWR _04511_ sky130_fd_sc_hd__nand2_1
X_17989_ clknet_leaf_8_clk _02273_ VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_127_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09412_ _04483_ _04812_ _04989_ CPU.cycles\[14\] VGND VGND VPWR VPWR _05115_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_140_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09343_ _05048_ VGND VGND VPWR VPWR _05049_ sky130_fd_sc_hd__buf_4
XFILLER_0_158_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_158_Right_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09274_ net1717 _04982_ _04983_ VGND VGND VPWR VPWR _04984_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14810__903 clknet_1_0__leaf__02696_ VGND VGND VPWR VPWR net935 sky130_fd_sc_hd__inv_2
XFILLER_0_7_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14203__380 clknet_1_0__leaf__08430_ VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__inv_2
XFILLER_0_105_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12750__203 clknet_1_1__leaf__07221_ VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__inv_2
X_08989_ CPU.aluReg\[29\] _04681_ _04706_ _04700_ VGND VGND VPWR VPWR _04707_ sky130_fd_sc_hd__a211o_1
X_10951_ net1545 _05733_ _06142_ VGND VGND VPWR VPWR _06176_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13670_ CPU.registerFile\[21\]\[23\] _07362_ _08089_ _07650_ VGND VGND VPWR VPWR
+ _08090_ sky130_fd_sc_hd__o22a_1
X_10882_ net2139 _05733_ _06105_ VGND VGND VPWR VPWR _06139_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__02696_ clknet_0__02696_ VGND VGND VPWR VPWR clknet_1_0__leaf__02696_
+ sky130_fd_sc_hd__clkbuf_16
X_12621_ _06515_ VGND VGND VPWR VPWR _07135_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_0__f__07223_ clknet_0__07223_ VGND VGND VPWR VPWR clknet_1_0__leaf__07223_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_66_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_125_Right_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15340_ CPU.registerFile\[20\]\[0\] CPU.registerFile\[21\]\[0\] _02829_ VGND VGND
+ VPWR VPWR _02839_ sky130_fd_sc_hd__mux2_1
X_12552_ net2436 _05026_ _07096_ VGND VGND VPWR VPWR _07099_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11503_ CPU.mem_rstrb _04689_ _06469_ VGND VGND VPWR VPWR _06470_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_136_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15271_ _02769_ VGND VGND VPWR VPWR _02770_ sky130_fd_sc_hd__buf_4
XFILLER_0_108_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12483_ _07062_ VGND VGND VPWR VPWR _01348_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17010_ net268 _01332_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_78_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11434_ _06432_ VGND VGND VPWR VPWR _06433_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_78_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14153_ _07127_ VGND VGND VPWR VPWR _08413_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11365_ _05737_ _06395_ VGND VGND VPWR VPWR _06396_ sky130_fd_sc_hd__nand2_2
X_13104_ CPU.registerFile\[1\]\[6\] _07256_ _07540_ _07258_ VGND VGND VPWR VPWR _07541_
+ sky130_fd_sc_hd__a22o_1
X_10316_ _05493_ net2323 _05777_ VGND VGND VPWR VPWR _05779_ sky130_fd_sc_hd__mux2_1
X_11296_ _05488_ _05738_ VGND VGND VPWR VPWR _06359_ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_91_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ _07359_ VGND VGND VPWR VPWR _07474_ sky130_fd_sc_hd__buf_4
X_17912_ net1101 _02196_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[30\] sky130_fd_sc_hd__dfxtp_1
X_10247_ _05493_ net1805 _05740_ VGND VGND VPWR VPWR _05742_ sky130_fd_sc_hd__mux2_1
X_17843_ net1032 _02127_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_10178_ net2450 _05694_ _05692_ VGND VGND VPWR VPWR _05695_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15192__105 clknet_1_0__leaf__02750_ VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__inv_2
X_17774_ net963 _02058_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16725_ _03995_ _05182_ _07132_ VGND VGND VPWR VPWR _04047_ sky130_fd_sc_hd__o21ai_1
X_13937_ CPU.registerFile\[31\]\[31\] _07502_ _07503_ CPU.registerFile\[27\]\[31\]
+ _07345_ VGND VGND VPWR VPWR _08349_ sky130_fd_sc_hd__o221a_1
XFILLER_0_135_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13868_ CPU.registerFile\[15\]\[29\] _07236_ _07239_ CPU.registerFile\[11\]\[29\]
+ _07820_ VGND VGND VPWR VPWR _08282_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_122_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12819_ net14 VGND VGND VPWR VPWR _07262_ sky130_fd_sc_hd__clkbuf_4
X_15607_ _03095_ _03099_ _02810_ VGND VGND VPWR VPWR _03100_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13799_ CPU.registerFile\[16\]\[27\] CPU.registerFile\[20\]\[27\] _07648_ VGND VGND
+ VPWR VPWR _08215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18326_ clknet_leaf_6_clk _02606_ VGND VGND VPWR VPWR per_uart.tx_busy sky130_fd_sc_hd__dfxtp_1
X_15538_ CPU.registerFile\[16\]\[4\] CPU.registerFile\[18\]\[4\] _03032_ VGND VGND
+ VPWR VPWR _03033_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15469_ _05093_ VGND VGND VPWR VPWR _02965_ sky130_fd_sc_hd__buf_4
X_18257_ net98 _02537_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17208_ net398 _01496_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_18188_ net219 _02468_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold603 CPU.registerFile\[3\]\[23\] VGND VGND VPWR VPWR net1844 sky130_fd_sc_hd__dlygate4sd3_1
X_17139_ net363 _01427_ VGND VGND VPWR VPWR CPU.aluReg\[3\] sky130_fd_sc_hd__dfxtp_1
Xhold614 CPU.registerFile\[26\]\[7\] VGND VGND VPWR VPWR net1855 sky130_fd_sc_hd__dlygate4sd3_1
Xhold625 CPU.registerFile\[26\]\[24\] VGND VGND VPWR VPWR net1866 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold636 CPU.registerFile\[31\]\[7\] VGND VGND VPWR VPWR net1877 sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 CPU.registerFile\[29\]\[13\] VGND VGND VPWR VPWR net1888 sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 CPU.registerFile\[27\]\[16\] VGND VGND VPWR VPWR net1899 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09961_ _05516_ net1838 _05570_ VGND VGND VPWR VPWR _05573_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold669 CPU.registerFile\[18\]\[6\] VGND VGND VPWR VPWR net1910 sky130_fd_sc_hd__dlygate4sd3_1
X_08912_ _04522_ _04534_ VGND VGND VPWR VPWR _04632_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09892_ _05529_ VGND VGND VPWR VPWR _02491_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__02659_ clknet_0__02659_ VGND VGND VPWR VPWR clknet_1_1__leaf__02659_
+ sky130_fd_sc_hd__clkbuf_16
X_14569__686 clknet_1_1__leaf__02672_ VGND VGND VPWR VPWR net718 sky130_fd_sc_hd__inv_2
X_08843_ CPU.aluIn1\[17\] _04494_ VGND VGND VPWR VPWR _04563_ sky130_fd_sc_hd__xnor2_1
Xhold1303 mapped_spi_flash.snd_bitcount\[0\] VGND VGND VPWR VPWR net2544 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08774_ CPU.Bimm\[12\] VGND VGND VPWR VPWR _04494_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_0_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780__229 clknet_1_1__leaf__07225_ VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09326_ _04250_ _04699_ _04808_ CPU.aluReg\[18\] _05032_ VGND VGND VPWR VPWR _05033_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14734__834 clknet_1_1__leaf__02689_ VGND VGND VPWR VPWR net866 sky130_fd_sc_hd__inv_2
XFILLER_0_63_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09257_ _04244_ _04210_ _04217_ CPU.aluReg\[21\] _04966_ VGND VGND VPWR VPWR _04967_
+ sky130_fd_sc_hd__a221o_1
Xclone36 _04655_ VGND VGND VPWR VPWR net1277 sky130_fd_sc_hd__buf_2
XFILLER_0_145_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_153_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09188_ CPU.PC\[16\] _04842_ VGND VGND VPWR VPWR _04900_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11150_ CPU.registerFile\[8\]\[4\] _05727_ _06274_ VGND VGND VPWR VPWR _06282_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10101_ CPU.registerFile\[18\]\[18\] _05046_ _05644_ VGND VGND VPWR VPWR _05648_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_73_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11081_ net1640 _05727_ _06237_ VGND VGND VPWR VPWR _06245_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10032_ net2157 _05046_ _05607_ VGND VGND VPWR VPWR _05611_ sky130_fd_sc_hd__mux2_1
X_14780__876 clknet_1_0__leaf__02693_ VGND VGND VPWR VPWR net908 sky130_fd_sc_hd__inv_2
X_14840_ clknet_1_0__leaf__02697_ VGND VGND VPWR VPWR _02700_ sky130_fd_sc_hd__buf_1
X_11983_ _05008_ net1703 _06758_ VGND VGND VPWR VPWR _06760_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13722_ _07394_ _08126_ _08140_ _08015_ VGND VGND VPWR VPWR _08141_ sky130_fd_sc_hd__a211o_1
X_10934_ _06167_ VGND VGND VPWR VPWR _02040_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_104_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17490_ net679 _01778_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__02748_ clknet_0__02748_ VGND VGND VPWR VPWR clknet_1_0__leaf__02748_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_104_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16441_ _08401_ _03906_ _03909_ _02934_ VGND VGND VPWR VPWR _03910_ sky130_fd_sc_hd__o211a_1
X_13653_ CPU.registerFile\[28\]\[22\] CPU.registerFile\[24\]\[22\] _07292_ VGND VGND
+ VPWR VPWR _08074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_27_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10865_ _06130_ VGND VGND VPWR VPWR _02072_ sky130_fd_sc_hd__clkbuf_1
X_14026__305 clknet_1_1__leaf__08362_ VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__inv_2
XFILLER_0_155_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__02679_ clknet_0__02679_ VGND VGND VPWR VPWR clknet_1_0__leaf__02679_
+ sky130_fd_sc_hd__clkbuf_16
X_12604_ _06577_ _07124_ _05942_ VGND VGND VPWR VPWR _00011_ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16372_ CPU.registerFile\[27\]\[28\] CPU.registerFile\[31\]\[28\] _08403_ VGND VGND
+ VPWR VPWR _03843_ sky130_fd_sc_hd__mux2_1
X_13584_ CPU.registerFile\[30\]\[20\] CPU.registerFile\[26\]\[20\] _07292_ VGND VGND
+ VPWR VPWR _08007_ sky130_fd_sc_hd__mux2_1
X_10796_ _05535_ CPU.registerFile\[30\]\[10\] _06092_ VGND VGND VPWR VPWR _06094_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15323_ _02813_ VGND VGND VPWR VPWR _02822_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18111_ net174 _02391_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_12535_ net2385 _04747_ _07085_ VGND VGND VPWR VPWR _07090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18042_ net1215 _02322_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_12466_ _07053_ VGND VGND VPWR VPWR _01356_ sky130_fd_sc_hd__clkbuf_1
X_15173__1199 clknet_1_1__leaf__02747_ VGND VGND VPWR VPWR net1231 sky130_fd_sc_hd__inv_2
XFILLER_0_2_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11417_ _05541_ net2465 _06419_ VGND VGND VPWR VPWR _06424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15185_ clknet_leaf_0_clk VGND VGND VPWR VPWR _02749_ sky130_fd_sc_hd__buf_1
X_12397_ _04731_ net2096 _07013_ VGND VGND VPWR VPWR _07017_ sky130_fd_sc_hd__mux2_1
X_14136_ _08399_ VGND VGND VPWR VPWR _08400_ sky130_fd_sc_hd__buf_4
X_11348_ _05541_ net2444 _06382_ VGND VGND VPWR VPWR _06387_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11279_ _06350_ VGND VGND VPWR VPWR _01878_ sky130_fd_sc_hd__clkbuf_1
X_15200__112 clknet_1_1__leaf__02751_ VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__inv_2
X_13018_ _07240_ VGND VGND VPWR VPWR _07457_ sky130_fd_sc_hd__clkbuf_8
X_17826_ net1015 _02110_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17757_ net946 _02041_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16708_ _03990_ VGND VGND VPWR VPWR _04032_ sky130_fd_sc_hd__buf_2
X_08490_ _04209_ VGND VGND VPWR VPWR _04210_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17688_ net877 _01976_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09111_ CPU.PC\[21\] _04822_ VGND VGND VPWR VPWR _04823_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18309_ clknet_leaf_16_clk _02589_ VGND VGND VPWR VPWR CPU.PC\[9\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_155_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09042_ _04232_ _04214_ _04754_ _04756_ VGND VGND VPWR VPWR _04757_ sky130_fd_sc_hd__a211o_1
XFILLER_0_143_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold400 CPU.registerFile\[4\]\[0\] VGND VGND VPWR VPWR net1641 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold411 CPU.registerFile\[6\]\[22\] VGND VGND VPWR VPWR net1652 sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 CPU.registerFile\[2\]\[26\] VGND VGND VPWR VPWR net1663 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold433 CPU.registerFile\[2\]\[29\] VGND VGND VPWR VPWR net1674 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 _02633_ VGND VGND VPWR VPWR net1685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 CPU.registerFile\[7\]\[5\] VGND VGND VPWR VPWR net1696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 CPU.registerFile\[10\]\[24\] VGND VGND VPWR VPWR net1707 sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 CPU.registerFile\[14\]\[21\] VGND VGND VPWR VPWR net1718 sky130_fd_sc_hd__dlygate4sd3_1
X_09944_ _05499_ net1831 _05559_ VGND VGND VPWR VPWR _05564_ sky130_fd_sc_hd__mux2_1
Xhold488 CPU.registerFile\[22\]\[20\] VGND VGND VPWR VPWR net1729 sky130_fd_sc_hd__dlygate4sd3_1
Xhold499 CPU.registerFile\[8\]\[27\] VGND VGND VPWR VPWR net1740 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09875_ _05045_ VGND VGND VPWR VPWR _05518_ sky130_fd_sc_hd__buf_6
Xhold1100 CPU.registerFile\[21\]\[7\] VGND VGND VPWR VPWR net2341 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1111 CPU.registerFile\[10\]\[13\] VGND VGND VPWR VPWR net2352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1122 CPU.registerFile\[21\]\[8\] VGND VGND VPWR VPWR net2363 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08826_ _04511_ _04545_ VGND VGND VPWR VPWR _04546_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_51_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1133 CPU.aluShamt\[2\] VGND VGND VPWR VPWR net2374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1144 CPU.registerFile\[4\]\[27\] VGND VGND VPWR VPWR net2385 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1155 CPU.registerFile\[21\]\[16\] VGND VGND VPWR VPWR net2396 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1166 CPU.registerFile\[25\]\[6\] VGND VGND VPWR VPWR net2407 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1177 CPU.registerFile\[10\]\[12\] VGND VGND VPWR VPWR net2418 sky130_fd_sc_hd__dlygate4sd3_1
X_08757_ _04380_ _04476_ _04226_ VGND VGND VPWR VPWR _04477_ sky130_fd_sc_hd__o21a_1
Xhold1188 CPU.registerFile\[25\]\[8\] VGND VGND VPWR VPWR net2429 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_306 _07418_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1199 CPU.registerFile\[15\]\[18\] VGND VGND VPWR VPWR net2440 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_317 _07914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_328 _08322_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_339 _03056_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08688_ net1292 CPU.aluIn1\[2\] VGND VGND VPWR VPWR _04408_ sky130_fd_sc_hd__and2b_1
XFILLER_0_95_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10650_ mapped_spi_flash.div_counter\[3\] mapped_spi_flash.div_counter\[2\] mapped_spi_flash.div_counter\[5\]
+ mapped_spi_flash.div_counter\[4\] VGND VGND VPWR VPWR _06010_ sky130_fd_sc_hd__or4_1
X_14322__463 clknet_1_0__leaf__08465_ VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__inv_2
XFILLER_0_64_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09309_ _04800_ _05014_ _05016_ _04768_ VGND VGND VPWR VPWR _05017_ sky130_fd_sc_hd__o211a_1
XFILLER_0_146_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10581_ net1316 _05970_ VGND VGND VPWR VPWR _05972_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13960__245 clknet_1_1__leaf__08356_ VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__inv_2
X_12320_ _06975_ VGND VGND VPWR VPWR _01424_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12251_ CPU.aluIn1\[16\] _06922_ _06894_ VGND VGND VPWR VPWR _06923_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11202_ _06309_ VGND VGND VPWR VPWR _01914_ sky130_fd_sc_hd__clkbuf_1
X_12182_ _04302_ _06865_ _06862_ _06869_ VGND VGND VPWR VPWR _01490_ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11133_ net2458 _05710_ _06263_ VGND VGND VPWR VPWR _06273_ sky130_fd_sc_hd__mux2_1
X_16990_ clknet_leaf_21_clk _01316_ VGND VGND VPWR VPWR CPU.rs2\[21\] sky130_fd_sc_hd__dfxtp_1
X_11064_ net2359 _05710_ _06226_ VGND VGND VPWR VPWR _06236_ sky130_fd_sc_hd__mux2_1
X_15941_ _05093_ _03422_ _03423_ _03424_ _03028_ VGND VGND VPWR VPWR _03425_ sky130_fd_sc_hd__o221a_1
X_10015_ net1870 _04762_ _05596_ VGND VGND VPWR VPWR _05602_ sky130_fd_sc_hd__mux2_1
X_15872_ CPU.registerFile\[16\]\[13\] _03068_ _03069_ CPU.registerFile\[17\]\[13\]
+ _02854_ VGND VGND VPWR VPWR _03358_ sky130_fd_sc_hd__o221a_1
X_17611_ net800 _01899_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12763__213 clknet_1_0__leaf__07224_ VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__inv_2
XFILLER_0_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17542_ net731 _01830_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_86_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11966_ _04731_ net2018 _06747_ VGND VGND VPWR VPWR _06751_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_86_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14405__538 clknet_1_1__leaf__02656_ VGND VGND VPWR VPWR net570 sky130_fd_sc_hd__inv_2
X_10917_ _06158_ VGND VGND VPWR VPWR _02048_ sky130_fd_sc_hd__clkbuf_1
X_13705_ _07650_ _08122_ _08123_ VGND VGND VPWR VPWR _08124_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_129_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17473_ net662 _01761_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[28\] sky130_fd_sc_hd__dfxtp_1
X_11897_ _06714_ VGND VGND VPWR VPWR _01621_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16424_ _02914_ _03891_ _03893_ _02864_ VGND VGND VPWR VPWR _03894_ sky130_fd_sc_hd__a211o_1
X_13636_ CPU.registerFile\[16\]\[22\] CPU.registerFile\[20\]\[22\] _07785_ VGND VGND
+ VPWR VPWR _08057_ sky130_fd_sc_hd__mux2_1
X_10848_ _06121_ VGND VGND VPWR VPWR _02080_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13567_ CPU.registerFile\[4\]\[20\] _07374_ VGND VGND VPWR VPWR _07990_ sky130_fd_sc_hd__or2_1
X_16355_ _03822_ _03826_ _02843_ VGND VGND VPWR VPWR _03827_ sky130_fd_sc_hd__a21o_1
X_14297__440 clknet_1_0__leaf__08463_ VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__inv_2
X_10779_ _05518_ net1655 _06081_ VGND VGND VPWR VPWR _06085_ sky130_fd_sc_hd__mux2_1
X_12518_ _07080_ VGND VGND VPWR VPWR _01331_ sky130_fd_sc_hd__clkbuf_1
X_15306_ net15 VGND VGND VPWR VPWR _02805_ sky130_fd_sc_hd__clkbuf_4
X_16286_ _02818_ _03758_ _03759_ VGND VGND VPWR VPWR _03760_ sky130_fd_sc_hd__a21o_1
XFILLER_0_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13498_ CPU.registerFile\[18\]\[18\] CPU.registerFile\[22\]\[18\] _07457_ VGND VGND
+ VPWR VPWR _07923_ sky130_fd_sc_hd__mux2_1
X_15129__1159 clknet_1_0__leaf__02743_ VGND VGND VPWR VPWR net1191 sky130_fd_sc_hd__inv_2
XFILLER_0_23_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18025_ net1198 _02305_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_12449_ _05381_ net1981 _07035_ VGND VGND VPWR VPWR _07044_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14119_ _08388_ VGND VGND VPWR VPWR _01468_ sky130_fd_sc_hd__clkbuf_1
X_15099_ _07188_ _02736_ _02727_ VGND VGND VPWR VPWR _02279_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_130_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14763__860 clknet_1_0__leaf__02692_ VGND VGND VPWR VPWR net892 sky130_fd_sc_hd__inv_2
X_09660_ _04419_ _05352_ VGND VGND VPWR VPWR _05353_ sky130_fd_sc_hd__xor2_1
X_08611_ CPU.aluIn1\[15\] _04255_ VGND VGND VPWR VPWR _04331_ sky130_fd_sc_hd__or2_1
X_16523__190 clknet_1_1__leaf__03964_ VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__inv_2
X_17809_ net998 _02093_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_09591_ net1274 _04292_ _04653_ VGND VGND VPWR VPWR _05286_ sky130_fd_sc_hd__nor3_2
X_08542_ CPU.aluIn1\[12\] _04261_ VGND VGND VPWR VPWR _04262_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08473_ _04194_ VGND VGND VPWR VPWR _02647_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_137_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_914 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_122_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09025_ _04358_ _04740_ VGND VGND VPWR VPWR _04741_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold230 _02168_ VGND VGND VPWR VPWR net1471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 mapped_spi_ram.rcv_data\[22\] VGND VGND VPWR VPWR net1482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 CPU.rs2\[30\] VGND VGND VPWR VPWR net1493 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 CPU.aluShamt\[0\] VGND VGND VPWR VPWR net1504 sky130_fd_sc_hd__dlygate4sd3_1
X_14846__935 clknet_1_0__leaf__02700_ VGND VGND VPWR VPWR net967 sky130_fd_sc_hd__inv_2
Xhold274 per_uart.uart0.rx_busy VGND VGND VPWR VPWR net1515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 CPU.rs2\[13\] VGND VGND VPWR VPWR net1526 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold296 _04111_ VGND VGND VPWR VPWR net1537 sky130_fd_sc_hd__dlygate4sd3_1
X_09927_ _05425_ VGND VGND VPWR VPWR _05553_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_148_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09858_ _05506_ VGND VGND VPWR VPWR _02502_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_29_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08809_ CPU.Iimm\[2\] CPU.Bimm\[2\] CPU.instr\[5\] VGND VGND VPWR VPWR _04529_ sky130_fd_sc_hd__mux2_4
XFILLER_0_99_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09789_ _05465_ VGND VGND VPWR VPWR _02530_ sky130_fd_sc_hd__clkbuf_1
X_15172__1198 clknet_1_1__leaf__02747_ VGND VGND VPWR VPWR net1230 sky130_fd_sc_hd__inv_2
X_11820_ _05448_ net1790 _06638_ VGND VGND VPWR VPWR _06673_ sky130_fd_sc_hd__mux2_1
XANTENNA_103 _05384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_114 _05448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_125 _05539_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_136 _05696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_147 _07260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_158 _07296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11751_ _06635_ _06636_ net2504 VGND VGND VPWR VPWR _06637_ sky130_fd_sc_hd__mux2_1
XANTENNA_169 _07398_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10702_ _05509_ net1813 _06034_ VGND VGND VPWR VPWR _06044_ sky130_fd_sc_hd__mux2_1
X_14892__977 clknet_1_0__leaf__02704_ VGND VGND VPWR VPWR net1009 sky130_fd_sc_hd__inv_2
XFILLER_0_154_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11682_ _06515_ VGND VGND VPWR VPWR _06594_ sky130_fd_sc_hd__buf_2
XFILLER_0_49_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13421_ CPU.registerFile\[14\]\[15\] CPU.registerFile\[10\]\[15\] _07274_ VGND VGND
+ VPWR VPWR _07849_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10633_ mapped_spi_flash.rcv_data\[7\] _05994_ VGND VGND VPWR VPWR _06001_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16140_ CPU.registerFile\[6\]\[21\] _03057_ _03140_ _03617_ VGND VGND VPWR VPWR _03618_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13352_ CPU.registerFile\[1\]\[13\] _07255_ _07781_ _07318_ VGND VGND VPWR VPWR _07782_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10564_ net1459 _05950_ _05952_ _05958_ VGND VGND VPWR VPWR _02200_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_101_Left_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12303_ net2517 _06962_ _06861_ VGND VGND VPWR VPWR _06963_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16071_ CPU.registerFile\[9\]\[19\] _08404_ _02860_ VGND VGND VPWR VPWR _03551_ sky130_fd_sc_hd__o21a_1
X_13283_ _07364_ _07714_ VGND VGND VPWR VPWR _07715_ sky130_fd_sc_hd__or2_1
X_10495_ CPU.aluIn1\[9\] CPU.Bimm\[9\] VGND VGND VPWR VPWR _05903_ sky130_fd_sc_hd__and2_1
X_12234_ CPU.aluReg\[21\] CPU.aluReg\[19\] _06906_ VGND VGND VPWR VPWR _06910_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12165_ _04284_ _06856_ VGND VGND VPWR VPWR _06857_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_112_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11116_ _06264_ VGND VGND VPWR VPWR _01955_ sky130_fd_sc_hd__clkbuf_1
X_12096_ _04659_ net2261 _06819_ VGND VGND VPWR VPWR _06820_ sky130_fd_sc_hd__mux2_1
X_16973_ clknet_leaf_26_clk _01299_ VGND VGND VPWR VPWR CPU.mem_wdata\[4\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_127_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15924_ CPU.registerFile\[1\]\[15\] _02867_ _03407_ _02895_ VGND VGND VPWR VPWR _03408_
+ sky130_fd_sc_hd__a22o_1
X_11047_ _06227_ VGND VGND VPWR VPWR _01987_ sky130_fd_sc_hd__clkbuf_1
X_15855_ _03336_ _03340_ _08410_ VGND VGND VPWR VPWR _03341_ sky130_fd_sc_hd__a21o_1
X_14806_ clknet_1_0__leaf__02686_ VGND VGND VPWR VPWR _02696_ sky130_fd_sc_hd__buf_1
X_15786_ CPU.registerFile\[30\]\[11\] CPU.registerFile\[26\]\[11\] _02787_ VGND VGND
+ VPWR VPWR _03274_ sky130_fd_sc_hd__mux2_1
X_12998_ CPU.registerFile\[7\]\[3\] _07262_ _07437_ _07265_ VGND VGND VPWR VPWR _07438_
+ sky130_fd_sc_hd__o211a_1
X_17525_ net714 _01813_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_11949_ _06741_ VGND VGND VPWR VPWR _01596_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17456_ net645 _01744_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16407_ _03252_ _03868_ _03876_ _02935_ VGND VGND VPWR VPWR _03877_ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13619_ CPU.registerFile\[5\]\[21\] CPU.registerFile\[4\]\[21\] _04986_ VGND VGND
+ VPWR VPWR _08041_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17387_ net576 _01675_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16338_ _02903_ _03799_ _03803_ _03809_ VGND VGND VPWR VPWR _03810_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16269_ CPU.registerFile\[29\]\[25\] _02772_ VGND VGND VPWR VPWR _03743_ sky130_fd_sc_hd__or2_1
X_14004__285 clknet_1_0__leaf__08360_ VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__inv_2
X_18008_ net1181 _02288_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09712_ net1630 _05402_ _05189_ VGND VGND VPWR VPWR _05403_ sky130_fd_sc_hd__mux2_1
X_09643_ mapped_spi_ram.rcv_data\[12\] net18 _04690_ mapped_spi_flash.rcv_data\[12\]
+ VGND VGND VPWR VPWR _05336_ sky130_fd_sc_hd__a22o_2
X_09574_ _04818_ _05257_ _05259_ _04955_ _05269_ VGND VGND VPWR VPWR _05270_ sky130_fd_sc_hd__o221a_1
XFILLER_0_78_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_143_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14927__1009 clknet_1_1__leaf__02707_ VGND VGND VPWR VPWR net1041 sky130_fd_sc_hd__inv_2
X_08525_ CPU.aluIn1\[21\] _04243_ VGND VGND VPWR VPWR _04245_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16600__70 clknet_1_1__leaf__03971_ VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__inv_2
XFILLER_0_34_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09008_ _04362_ _04230_ _04360_ VGND VGND VPWR VPWR _04725_ sky130_fd_sc_hd__or3_1
XFILLER_0_130_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10280_ _05526_ net1766 _05751_ VGND VGND VPWR VPWR _05759_ sky130_fd_sc_hd__mux2_1
X_14434__564 clknet_1_0__leaf__02659_ VGND VGND VPWR VPWR net596 sky130_fd_sc_hd__inv_2
XFILLER_0_130_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12921_ _07361_ VGND VGND VPWR VPWR _07362_ sky130_fd_sc_hd__buf_4
X_15128__1158 clknet_1_0__leaf__02743_ VGND VGND VPWR VPWR net1190 sky130_fd_sc_hd__inv_2
X_15640_ CPU.registerFile\[24\]\[7\] _03130_ _02790_ _03131_ VGND VGND VPWR VPWR _03132_
+ sky130_fd_sc_hd__o211a_1
X_12852_ CPU.registerFile\[31\]\[0\] _07289_ _07290_ CPU.registerFile\[27\]\[0\] _07294_
+ VGND VGND VPWR VPWR _07295_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_83_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14900__984 clknet_1_1__leaf__02705_ VGND VGND VPWR VPWR net1016 sky130_fd_sc_hd__inv_2
X_11803_ _06664_ VGND VGND VPWR VPWR _01665_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15571_ _03064_ VGND VGND VPWR VPWR _03065_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17310_ net499 _01598_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11734_ mapped_spi_ram.state\[3\] _06472_ _06569_ VGND VGND VPWR VPWR _06625_ sky130_fd_sc_hd__o21a_1
XFILLER_0_84_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18290_ net123 _02570_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17241_ net431 _01529_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_11665_ mapped_spi_ram.rcv_data\[26\] _06577_ VGND VGND VPWR VPWR _06584_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13404_ _07271_ _07822_ _07825_ _07832_ _07766_ VGND VGND VPWR VPWR _07833_ sky130_fd_sc_hd__o311a_1
X_10616_ mapped_spi_flash.rcv_data\[14\] _05981_ VGND VGND VPWR VPWR _05991_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17172_ clknet_leaf_24_clk _01460_ VGND VGND VPWR VPWR CPU.instr\[2\] sky130_fd_sc_hd__dfxtp_2
X_11596_ net1381 _06517_ _06508_ _06535_ VGND VGND VPWR VPWR _06536_ sky130_fd_sc_hd__a211o_1
X_14517__639 clknet_1_0__leaf__02667_ VGND VGND VPWR VPWR net671 sky130_fd_sc_hd__inv_2
XFILLER_0_91_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16123_ CPU.registerFile\[8\]\[21\] _02789_ _03117_ _03600_ VGND VGND VPWR VPWR _03601_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13335_ _07305_ VGND VGND VPWR VPWR _07766_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10547_ mapped_spi_flash.snd_bitcount\[4\] _05944_ VGND VGND VPWR VPWR _05945_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_114_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14255__427 clknet_1_0__leaf__08435_ VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__inv_2
X_16054_ CPU.registerFile\[7\]\[19\] _02898_ _02887_ _03533_ VGND VGND VPWR VPWR _03534_
+ sky130_fd_sc_hd__o211a_1
X_13266_ CPU.registerFile\[14\]\[10\] CPU.registerFile\[10\]\[10\] _07492_ VGND VGND
+ VPWR VPWR _07699_ sky130_fd_sc_hd__mux2_1
X_10478_ CPU.PC\[12\] _05867_ _05888_ _04551_ VGND VGND VPWR VPWR _05889_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_110_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__02692_ clknet_0__02692_ VGND VGND VPWR VPWR clknet_1_1__leaf__02692_
+ sky130_fd_sc_hd__clkbuf_16
X_12217_ CPU.aluReg\[25\] CPU.aluReg\[23\] _06871_ VGND VGND VPWR VPWR _06897_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_94_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13197_ CPU.registerFile\[30\]\[8\] CPU.registerFile\[26\]\[8\] _07492_ VGND VGND
+ VPWR VPWR _07632_ sky130_fd_sc_hd__mux2_1
X_12148_ _05306_ net1938 _06841_ VGND VGND VPWR VPWR _06847_ sky130_fd_sc_hd__mux2_1
X_16956_ net251 _01282_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[19\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12079_ _06810_ VGND VGND VPWR VPWR _01534_ sky130_fd_sc_hd__clkbuf_1
X_15907_ _03065_ _03390_ _03391_ VGND VGND VPWR VPWR _03392_ sky130_fd_sc_hd__o21a_1
X_16887_ _04165_ _04164_ per_uart.uart0.rx_bitcount\[1\] per_uart.uart0.rx_bitcount\[0\]
+ VGND VGND VPWR VPWR _04168_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_139_Right_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15838_ CPU.registerFile\[16\]\[12\] _03068_ _03069_ CPU.registerFile\[17\]\[12\]
+ _02779_ VGND VGND VPWR VPWR _03325_ sky130_fd_sc_hd__o221a_1
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15769_ _03015_ _03255_ _03256_ _03257_ _02930_ VGND VGND VPWR VPWR _03258_ sky130_fd_sc_hd__a221o_1
X_14875__961 clknet_1_0__leaf__02703_ VGND VGND VPWR VPWR net993 sky130_fd_sc_hd__inv_2
X_17508_ net697 _01796_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_09290_ _04343_ _04488_ _04998_ _04768_ VGND VGND VPWR VPWR _04999_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16586__58 clknet_1_1__leaf__03969_ VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__inv_2
XFILLER_0_157_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_14 _02867_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17439_ net628 _01727_ VGND VGND VPWR VPWR mapped_spi_ram.snd_bitcount\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_25 _02948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_36 _03283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_47 _04730_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_880 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_58 _04981_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_69 _05108_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15171__1197 clknet_1_1__leaf__02747_ VGND VGND VPWR VPWR net1229 sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__08466_ clknet_0__08466_ VGND VGND VPWR VPWR clknet_1_1__leaf__08466_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_63_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_145_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_106_Right_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap16 _05068_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
X_09626_ _04800_ _05319_ VGND VGND VPWR VPWR _05320_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_39_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09557_ net2106 _05253_ _05189_ VGND VGND VPWR VPWR _05254_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08508_ CPU.aluIn1\[28\] _04227_ VGND VGND VPWR VPWR _04228_ sky130_fd_sc_hd__and2_1
X_09488_ _05187_ VGND VGND VPWR VPWR _05188_ sky130_fd_sc_hd__buf_4
XFILLER_0_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11450_ _06441_ VGND VGND VPWR VPWR _01798_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10401_ _04192_ VGND VGND VPWR VPWR _05830_ sky130_fd_sc_hd__buf_2
XFILLER_0_34_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11381_ _05505_ net2482 _06397_ VGND VGND VPWR VPWR _06405_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13120_ _07237_ VGND VGND VPWR VPWR _07557_ sky130_fd_sc_hd__buf_4
X_10332_ _05509_ net2246 _05777_ VGND VGND VPWR VPWR _05787_ sky130_fd_sc_hd__mux2_1
X_13051_ CPU.registerFile\[13\]\[4\] _07414_ _07488_ CPU.registerFile\[9\]\[4\] _07489_
+ VGND VGND VPWR VPWR _07490_ sky130_fd_sc_hd__o221a_1
X_10263_ _05509_ net1666 _05740_ VGND VGND VPWR VPWR _05750_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12002_ _05188_ net1726 _06769_ VGND VGND VPWR VPWR _06770_ sky130_fd_sc_hd__mux2_1
X_10194_ _05705_ VGND VGND VPWR VPWR _02333_ sky130_fd_sc_hd__clkbuf_1
X_16810_ _07178_ _08355_ net1529 VGND VGND VPWR VPWR _04116_ sky130_fd_sc_hd__o21ai_1
X_17790_ net979 _02074_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_14705__809 clknet_1_0__leaf__02685_ VGND VGND VPWR VPWR net841 sky130_fd_sc_hd__inv_2
XFILLER_0_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16741_ _04056_ _04060_ _04015_ VGND VGND VPWR VPWR _02593_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12904_ CPU.registerFile\[31\]\[1\] _07289_ _07290_ CPU.registerFile\[27\]\[1\] _07345_
+ VGND VGND VPWR VPWR _07346_ sky130_fd_sc_hd__o221a_1
X_16672_ _04001_ _05369_ _03990_ VGND VGND VPWR VPWR _04002_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13884_ _07322_ _08296_ VGND VGND VPWR VPWR _08297_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15623_ CPU.aluIn1\[6\] _03081_ _03115_ _03080_ VGND VGND VPWR VPWR _02420_ sky130_fd_sc_hd__o211a_1
X_12835_ _07252_ VGND VGND VPWR VPWR _07278_ sky130_fd_sc_hd__buf_4
XFILLER_0_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_26_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_8
X_18342_ clknet_leaf_5_clk _02622_ VGND VGND VPWR VPWR per_uart.rx_data\[6\] sky130_fd_sc_hd__dfxtp_1
X_15554_ CPU.registerFile\[24\]\[5\] _02789_ _02790_ _03047_ VGND VGND VPWR VPWR _03048_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11717_ mapped_spi_ram.rcv_data\[3\] _06601_ VGND VGND VPWR VPWR _06613_ sky130_fd_sc_hd__or2_1
X_18273_ net106 _02553_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_12697_ per_uart.uart0.tx_bitcount\[2\] per_uart.uart0.tx_bitcount\[1\] per_uart.uart0.tx_bitcount\[0\]
+ per_uart.uart0.tx_bitcount\[3\] VGND VGND VPWR VPWR _07179_ sky130_fd_sc_hd__and4bb_1
X_15485_ CPU.registerFile\[2\]\[3\] _02872_ _02980_ CPU.registerFile\[3\]\[3\] _02940_
+ VGND VGND VPWR VPWR _02981_ sky130_fd_sc_hd__a221o_1
XFILLER_0_126_223 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17224_ net414 _01512_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[17\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_0__03962_ _03962_ VGND VGND VPWR VPWR clknet_0__03962_ sky130_fd_sc_hd__clkbuf_16
X_11648_ mapped_spi_ram.rcv_bitcount\[5\] mapped_spi_ram.rcv_bitcount\[4\] _06571_
+ VGND VGND VPWR VPWR _06572_ sky130_fd_sc_hd__or3_1
XFILLER_0_141_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17155_ net379 _01443_ VGND VGND VPWR VPWR CPU.aluReg\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_96_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11579_ _06494_ VGND VGND VPWR VPWR _06524_ sky130_fd_sc_hd__buf_2
XFILLER_0_3_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold807 CPU.registerFile\[12\]\[19\] VGND VGND VPWR VPWR net2048 sky130_fd_sc_hd__dlygate4sd3_1
X_16106_ CPU.registerFile\[9\]\[20\] _08404_ _02860_ VGND VGND VPWR VPWR _03585_ sky130_fd_sc_hd__o21a_1
X_13318_ CPU.registerFile\[7\]\[12\] _07262_ _07748_ _05284_ VGND VGND VPWR VPWR _07749_
+ sky130_fd_sc_hd__o211a_1
Xhold818 CPU.registerFile\[15\]\[3\] VGND VGND VPWR VPWR net2059 sky130_fd_sc_hd__dlygate4sd3_1
Xhold829 CPU.registerFile\[2\]\[5\] VGND VGND VPWR VPWR net2070 sky130_fd_sc_hd__dlygate4sd3_1
X_17086_ net344 _01408_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[16\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__02744_ clknet_0__02744_ VGND VGND VPWR VPWR clknet_1_1__leaf__02744_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_40_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16037_ CPU.registerFile\[2\]\[18\] _03143_ _02980_ CPU.registerFile\[3\]\[18\] _03144_
+ VGND VGND VPWR VPWR _03518_ sky130_fd_sc_hd__a221o_1
X_14926__1008 clknet_1_0__leaf__02707_ VGND VGND VPWR VPWR net1040 sky130_fd_sc_hd__inv_2
X_13249_ CPU.registerFile\[23\]\[10\] _07382_ _07681_ _07418_ _07288_ VGND VGND VPWR
+ VPWR _07682_ sky130_fd_sc_hd__o221a_1
XFILLER_0_149_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__02675_ clknet_0__02675_ VGND VGND VPWR VPWR clknet_1_1__leaf__02675_
+ sky130_fd_sc_hd__clkbuf_16
X_08790_ CPU.aluIn1\[11\] CPU.Bimm\[12\] VGND VGND VPWR VPWR _04510_ sky130_fd_sc_hd__nand2_1
X_17988_ clknet_leaf_7_clk _02272_ VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_127_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16939_ net234 _01265_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_09411_ _04716_ _05113_ _04717_ VGND VGND VPWR VPWR _05114_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_140_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463__590 clknet_1_0__leaf__02662_ VGND VGND VPWR VPWR net622 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_140_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_17_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_94_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09342_ mapped_spi_ram.rcv_data\[9\] net18 _04690_ mapped_spi_flash.rcv_data\[9\]
+ VGND VGND VPWR VPWR _05048_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_48_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09273_ _04667_ VGND VGND VPWR VPWR _04983_ sky130_fd_sc_hd__buf_4
XFILLER_0_63_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14238__411 clknet_1_0__leaf__08434_ VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__inv_2
X_15127__1157 clknet_1_0__leaf__02743_ VGND VGND VPWR VPWR net1189 sky130_fd_sc_hd__inv_2
XFILLER_0_31_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08988_ _04226_ _04701_ _04705_ _04678_ VGND VGND VPWR VPWR _04706_ sky130_fd_sc_hd__a2bb2o_1
X_14546__665 clknet_1_1__leaf__02670_ VGND VGND VPWR VPWR net697 sky130_fd_sc_hd__inv_2
X_10950_ _06175_ VGND VGND VPWR VPWR _02032_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_3_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09609_ _05300_ _05301_ _05303_ _04708_ VGND VGND VPWR VPWR _05304_ sky130_fd_sc_hd__o31a_1
X_10881_ _06138_ VGND VGND VPWR VPWR _02064_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__02695_ clknet_0__02695_ VGND VGND VPWR VPWR clknet_1_0__leaf__02695_
+ sky130_fd_sc_hd__clkbuf_16
X_12620_ _04294_ _04830_ VGND VGND VPWR VPWR _07134_ sky130_fd_sc_hd__nand2_1
Xclkbuf_1_0__f__07222_ clknet_0__07222_ VGND VGND VPWR VPWR clknet_1_0__leaf__07222_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_155_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12551_ _07098_ VGND VGND VPWR VPWR _01283_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15078__1142 clknet_1_0__leaf__02724_ VGND VGND VPWR VPWR net1174 sky130_fd_sc_hd__inv_2
X_11502_ mapped_spi_ram.state\[2\] VGND VGND VPWR VPWR _06469_ sky130_fd_sc_hd__inv_2
X_16565__39 clknet_1_0__leaf__03967_ VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__inv_2
XFILLER_0_81_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12482_ net2184 _05694_ _07060_ VGND VGND VPWR VPWR _07062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15270_ _05439_ VGND VGND VPWR VPWR _02769_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_136_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11433_ _05775_ _06395_ VGND VGND VPWR VPWR _06432_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_78_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14711__813 clknet_1_0__leaf__02687_ VGND VGND VPWR VPWR net845 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_78_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14152_ _08412_ VGND VGND VPWR VPWR _01477_ sky130_fd_sc_hd__clkbuf_1
X_11364_ _04664_ CPU.writeBack _04665_ _04663_ VGND VGND VPWR VPWR _06395_ sky130_fd_sc_hd__and4b_2
X_14291__435 clknet_1_1__leaf__08462_ VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__inv_2
XFILLER_0_22_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13103_ CPU.registerFile\[5\]\[6\] CPU.registerFile\[4\]\[6\] _04986_ VGND VGND VPWR
+ VPWR _07540_ sky130_fd_sc_hd__mux2_1
X_10315_ _05778_ VGND VGND VPWR VPWR _02270_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11295_ _06358_ VGND VGND VPWR VPWR _01870_ sky130_fd_sc_hd__clkbuf_1
X_13034_ _07465_ _07472_ _07395_ VGND VGND VPWR VPWR _07473_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_91_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17911_ net1100 _02195_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[29\] sky130_fd_sc_hd__dfxtp_1
X_10246_ _05741_ VGND VGND VPWR VPWR _02317_ sky130_fd_sc_hd__clkbuf_1
X_17842_ net1031 _02126_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_10177_ _05007_ VGND VGND VPWR VPWR _05694_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_109_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17773_ net962 _02057_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16724_ _08379_ _05177_ _04006_ VGND VGND VPWR VPWR _04046_ sky130_fd_sc_hd__or3b_1
X_13936_ CPU.registerFile\[29\]\[31\] _07482_ _07420_ CPU.registerFile\[25\]\[31\]
+ _08347_ VGND VGND VPWR VPWR _08348_ sky130_fd_sc_hd__o221a_1
XFILLER_0_44_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15170__1196 clknet_1_0__leaf__02747_ VGND VGND VPWR VPWR net1228 sky130_fd_sc_hd__inv_2
X_13867_ CPU.registerFile\[14\]\[29\] CPU.registerFile\[10\]\[29\] _07480_ VGND VGND
+ VPWR VPWR _08281_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_122_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15606_ _02797_ _03096_ _03097_ _03098_ _03054_ VGND VGND VPWR VPWR _03099_ sky130_fd_sc_hd__a221o_1
X_12818_ CPU.registerFile\[2\]\[0\] CPU.registerFile\[3\]\[0\] _07260_ VGND VGND VPWR
+ VPWR _07261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13798_ CPU.registerFile\[23\]\[27\] _07282_ _08213_ VGND VGND VPWR VPWR _08214_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18325_ clknet_leaf_7_clk net1512 VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dfxtp_1
X_15537_ _05440_ VGND VGND VPWR VPWR _03032_ sky130_fd_sc_hd__buf_4
XFILLER_0_155_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18256_ net97 _02536_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_15468_ CPU.registerFile\[9\]\[3\] CPU.registerFile\[13\]\[3\] _02887_ VGND VGND
+ VPWR VPWR _02964_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17207_ net397 _01495_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_18187_ net218 _02467_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_15399_ CPU.registerFile\[20\]\[1\] CPU.registerFile\[22\]\[1\] _05440_ VGND VGND
+ VPWR VPWR _02897_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17138_ net362 _01426_ VGND VGND VPWR VPWR CPU.aluReg\[2\] sky130_fd_sc_hd__dfxtp_1
Xhold604 CPU.registerFile\[7\]\[29\] VGND VGND VPWR VPWR net1845 sky130_fd_sc_hd__dlygate4sd3_1
Xhold615 CPU.registerFile\[24\]\[30\] VGND VGND VPWR VPWR net1856 sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 CPU.registerFile\[3\]\[6\] VGND VGND VPWR VPWR net1867 sky130_fd_sc_hd__dlygate4sd3_1
Xhold637 CPU.registerFile\[7\]\[28\] VGND VGND VPWR VPWR net1878 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold648 CPU.registerFile\[24\]\[26\] VGND VGND VPWR VPWR net1889 sky130_fd_sc_hd__dlygate4sd3_1
X_09960_ _05572_ VGND VGND VPWR VPWR _02466_ sky130_fd_sc_hd__clkbuf_1
X_17069_ net327 _01391_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold659 CPU.registerFile\[17\]\[7\] VGND VGND VPWR VPWR net1900 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_6_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_8
X_08911_ CPU.PC\[3\] _04598_ _04628_ _04630_ VGND VGND VPWR VPWR _04631_ sky130_fd_sc_hd__o2bb2a_1
X_09891_ _05528_ net2324 _05512_ VGND VGND VPWR VPWR _05529_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__02658_ clknet_0__02658_ VGND VGND VPWR VPWR clknet_1_1__leaf__02658_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_139_Left_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08842_ _04558_ _04561_ VGND VGND VPWR VPWR _04562_ sky130_fd_sc_hd__nand2_2
Xclkbuf_0__02689_ _02689_ VGND VGND VPWR VPWR clknet_0__02689_ sky130_fd_sc_hd__clkbuf_16
X_08773_ _04212_ _04220_ _04490_ _04492_ VGND VGND VPWR VPWR _04493_ sky130_fd_sc_hd__o31a_1
XFILLER_0_26_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09325_ _04337_ _04683_ VGND VGND VPWR VPWR _05032_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09256_ _04450_ _04701_ VGND VGND VPWR VPWR _04966_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclone37 _04642_ VGND VGND VPWR VPWR net1290 sky130_fd_sc_hd__buf_2
X_09187_ _04845_ _04897_ _04898_ VGND VGND VPWR VPWR _04899_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_153_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10100_ _05647_ VGND VGND VPWR VPWR _02369_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_73_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11080_ _06244_ VGND VGND VPWR VPWR _01971_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_73_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10031_ _05610_ VGND VGND VPWR VPWR _02401_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11982_ _06759_ VGND VGND VPWR VPWR _01581_ sky130_fd_sc_hd__clkbuf_1
X_13721_ _07334_ _08129_ _08132_ _08139_ _07766_ VGND VGND VPWR VPWR _08140_ sky130_fd_sc_hd__o311a_1
X_10933_ net1547 _05715_ _06165_ VGND VGND VPWR VPWR _06167_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__02747_ clknet_0__02747_ VGND VGND VPWR VPWR clknet_1_0__leaf__02747_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_104_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16440_ _08405_ _03907_ _03908_ VGND VGND VPWR VPWR _03909_ sky130_fd_sc_hd__a21o_1
X_10864_ net2266 _05715_ _06128_ VGND VGND VPWR VPWR _06130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13652_ CPU.registerFile\[31\]\[22\] _07556_ _07557_ CPU.registerFile\[27\]\[22\]
+ _07345_ VGND VGND VPWR VPWR _08073_ sky130_fd_sc_hd__o221a_1
X_14925__1007 clknet_1_0__leaf__02707_ VGND VGND VPWR VPWR net1039 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_27_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__02678_ clknet_0__02678_ VGND VGND VPWR VPWR clknet_1_0__leaf__02678_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_156_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12603_ _06483_ mapped_spi_ram.state\[3\] _06499_ net1335 VGND VGND VPWR VPWR _07124_
+ sky130_fd_sc_hd__a22o_1
X_16371_ _02911_ _03839_ _03841_ _03245_ VGND VGND VPWR VPWR _03842_ sky130_fd_sc_hd__a211o_1
XFILLER_0_155_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13583_ CPU.registerFile\[13\]\[20\] _07282_ _08005_ VGND VGND VPWR VPWR _08006_
+ sky130_fd_sc_hd__o21a_1
X_10795_ _06093_ VGND VGND VPWR VPWR _02105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18110_ net173 _02390_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_15322_ _08394_ _05405_ VGND VGND VPWR VPWR _02821_ sky130_fd_sc_hd__nor2_4
X_12534_ _07089_ VGND VGND VPWR VPWR _01291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18041_ net1214 _02321_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_12465_ net2230 _05677_ _07049_ VGND VGND VPWR VPWR _07053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11416_ _06423_ VGND VGND VPWR VPWR _01814_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12396_ _07016_ VGND VGND VPWR VPWR _01389_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11347_ _06386_ VGND VGND VPWR VPWR _01846_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14135_ _05440_ VGND VGND VPWR VPWR _08399_ sky130_fd_sc_hd__clkbuf_4
X_11278_ CPU.registerFile\[9\]\[8\] _05719_ _06346_ VGND VGND VPWR VPWR _06350_ sky130_fd_sc_hd__mux2_1
X_10229_ _05380_ VGND VGND VPWR VPWR _05729_ sky130_fd_sc_hd__clkbuf_4
X_13017_ CPU.mem_wdata\[3\] _07229_ _07456_ _07135_ VGND VGND VPWR VPWR _01298_ sky130_fd_sc_hd__o211a_1
X_17825_ net1014 _02109_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_17756_ net945 _02040_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16707_ _04026_ _04031_ _04015_ VGND VGND VPWR VPWR _02588_ sky130_fd_sc_hd__a21oi_1
X_13919_ CPU.registerFile\[1\]\[31\] _07576_ _08330_ _07288_ VGND VGND VPWR VPWR _08331_
+ sky130_fd_sc_hd__a211o_1
X_17687_ net876 _01975_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_15126__1156 clknet_1_0__leaf__02743_ VGND VGND VPWR VPWR net1188 sky130_fd_sc_hd__inv_2
XFILLER_0_58_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09110_ CPU.Iimm\[1\] _04496_ _04820_ VGND VGND VPWR VPWR _04822_ sky130_fd_sc_hd__mux2_1
X_18308_ clknet_leaf_15_clk _02588_ VGND VGND VPWR VPWR CPU.PC\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_40_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09041_ _04355_ _04210_ _04218_ CPU.aluReg\[26\] _04755_ VGND VGND VPWR VPWR _04756_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_143_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18239_ net80 _02519_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14575__691 clknet_1_0__leaf__02673_ VGND VGND VPWR VPWR net723 sky130_fd_sc_hd__inv_2
XFILLER_0_72_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold401 CPU.registerFile\[26\]\[31\] VGND VGND VPWR VPWR net1642 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold412 CPU.registerFile\[28\]\[0\] VGND VGND VPWR VPWR net1653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold423 CPU.registerFile\[18\]\[30\] VGND VGND VPWR VPWR net1664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 CPU.registerFile\[5\]\[16\] VGND VGND VPWR VPWR net1675 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold445 CPU.registerFile\[16\]\[28\] VGND VGND VPWR VPWR net1686 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold456 CPU.registerFile\[30\]\[2\] VGND VGND VPWR VPWR net1697 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_147_Left_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold467 CPU.registerFile\[30\]\[15\] VGND VGND VPWR VPWR net1708 sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 CPU.registerFile\[16\]\[20\] VGND VGND VPWR VPWR net1719 sky130_fd_sc_hd__dlygate4sd3_1
X_09943_ _05563_ VGND VGND VPWR VPWR _02474_ sky130_fd_sc_hd__clkbuf_1
Xhold489 CPU.registerFile\[26\]\[20\] VGND VGND VPWR VPWR net1730 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09874_ _05517_ VGND VGND VPWR VPWR _02497_ sky130_fd_sc_hd__clkbuf_1
X_15077__1141 clknet_1_0__leaf__02724_ VGND VGND VPWR VPWR net1173 sky130_fd_sc_hd__inv_2
Xhold1101 CPU.registerFile\[28\]\[7\] VGND VGND VPWR VPWR net2342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1112 CPU.registerFile\[20\]\[23\] VGND VGND VPWR VPWR net2353 sky130_fd_sc_hd__dlygate4sd3_1
X_08825_ CPU.aluIn1\[10\] CPU.Bimm\[10\] VGND VGND VPWR VPWR _04545_ sky130_fd_sc_hd__or2_1
Xhold1123 CPU.registerFile\[17\]\[10\] VGND VGND VPWR VPWR net2364 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1134 CPU.registerFile\[23\]\[8\] VGND VGND VPWR VPWR net2375 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1145 CPU.registerFile\[17\]\[17\] VGND VGND VPWR VPWR net2386 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1156 CPU.registerFile\[18\]\[24\] VGND VGND VPWR VPWR net2397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1167 CPU.registerFile\[24\]\[19\] VGND VGND VPWR VPWR net2408 sky130_fd_sc_hd__dlygate4sd3_1
X_08756_ _04467_ _04475_ _04362_ VGND VGND VPWR VPWR _04476_ sky130_fd_sc_hd__a21oi_2
Xhold1178 CPU.registerFile\[31\]\[13\] VGND VGND VPWR VPWR net2419 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1189 CPU.registerFile\[25\]\[13\] VGND VGND VPWR VPWR net2430 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_307 _07418_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_318 _07914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_329 _08322_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08687_ _04286_ CPU.aluIn1\[3\] VGND VGND VPWR VPWR _04407_ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_156_Left_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14658__766 clknet_1_1__leaf__02681_ VGND VGND VPWR VPWR net798 sky130_fd_sc_hd__inv_2
XFILLER_0_153_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09308_ _04800_ _05015_ VGND VGND VPWR VPWR _05016_ sky130_fd_sc_hd__nand2_1
X_10580_ net1316 _05968_ _05971_ _05936_ VGND VGND VPWR VPWR _02197_ sky130_fd_sc_hd__o211a_1
X_09239_ _04943_ _04949_ _04773_ VGND VGND VPWR VPWR _04950_ sky130_fd_sc_hd__o21a_1
XFILLER_0_23_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12250_ CPU.aluReg\[17\] CPU.aluReg\[15\] _06906_ VGND VGND VPWR VPWR _06922_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11201_ _05530_ CPU.registerFile\[22\]\[12\] _06299_ VGND VGND VPWR VPWR _06309_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12181_ net1504 VGND VGND VPWR VPWR _06869_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11132_ _06272_ VGND VGND VPWR VPWR _01947_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold990 CPU.registerFile\[31\]\[19\] VGND VGND VPWR VPWR net2231 sky130_fd_sc_hd__dlygate4sd3_1
X_11063_ _06235_ VGND VGND VPWR VPWR _01979_ sky130_fd_sc_hd__clkbuf_1
X_15940_ CPU.registerFile\[20\]\[15\] _03025_ _02829_ VGND VGND VPWR VPWR _03424_
+ sky130_fd_sc_hd__a21o_1
X_14823__914 clknet_1_0__leaf__02698_ VGND VGND VPWR VPWR net946 sky130_fd_sc_hd__inv_2
X_10014_ _05601_ VGND VGND VPWR VPWR _02409_ sky130_fd_sc_hd__clkbuf_1
X_15871_ CPU.registerFile\[20\]\[13\] CPU.registerFile\[21\]\[13\] _03066_ VGND VGND
+ VPWR VPWR _03357_ sky130_fd_sc_hd__mux2_1
X_17610_ net799 _01898_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17541_ net730 _01829_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11965_ _06750_ VGND VGND VPWR VPWR _01589_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_86_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_86_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13704_ CPU.registerFile\[21\]\[24\] _07244_ _07429_ CPU.registerFile\[17\]\[24\]
+ _07349_ VGND VGND VPWR VPWR _08123_ sky130_fd_sc_hd__o221a_1
X_10916_ net1574 _05698_ _06154_ VGND VGND VPWR VPWR _06158_ sky130_fd_sc_hd__mux2_1
X_17472_ net661 _01760_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[27\] sky130_fd_sc_hd__dfxtp_1
X_14684_ clknet_1_1__leaf__02675_ VGND VGND VPWR VPWR _02684_ sky130_fd_sc_hd__buf_1
X_11896_ net2437 _05675_ _06711_ VGND VGND VPWR VPWR _06714_ sky130_fd_sc_hd__mux2_1
X_16423_ CPU.registerFile\[30\]\[29\] _05050_ _02923_ _03892_ VGND VGND VPWR VPWR
+ _03893_ sky130_fd_sc_hd__o211a_1
X_13635_ CPU.registerFile\[1\]\[22\] _07387_ _08055_ _07379_ VGND VGND VPWR VPWR _08056_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10847_ net2393 _05698_ _06117_ VGND VGND VPWR VPWR _06121_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16354_ _02770_ _03823_ _03824_ _03825_ _05093_ VGND VGND VPWR VPWR _03826_ sky130_fd_sc_hd__a221o_1
XFILLER_0_137_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13566_ _07801_ _07985_ _07986_ _07988_ _07555_ VGND VGND VPWR VPWR _07989_ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10778_ _06084_ VGND VGND VPWR VPWR _02113_ sky130_fd_sc_hd__clkbuf_1
X_15305_ CPU.registerFile\[25\]\[0\] _02802_ _02803_ VGND VGND VPWR VPWR _02804_ sky130_fd_sc_hd__o21a_1
X_12517_ net1783 _05729_ _07071_ VGND VGND VPWR VPWR _07080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16285_ CPU.registerFile\[2\]\[25\] _02821_ _02822_ CPU.registerFile\[3\]\[25\] _02874_
+ VGND VGND VPWR VPWR _03759_ sky130_fd_sc_hd__a221o_1
X_13497_ CPU.rs2\[17\] _07705_ _07907_ _07922_ _07737_ VGND VGND VPWR VPWR _01312_
+ sky130_fd_sc_hd__o221a_1
X_18024_ net1197 _02304_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_12448_ _07043_ VGND VGND VPWR VPWR _01364_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_117_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12379_ _05359_ net2158 _06999_ VGND VGND VPWR VPWR _07007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14118_ _04663_ _05191_ _08387_ VGND VGND VPWR VPWR _08388_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15098_ net1348 _07187_ VGND VGND VPWR VPWR _02736_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_130_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08610_ _04258_ _04328_ _04329_ VGND VGND VPWR VPWR _04330_ sky130_fd_sc_hd__a21boi_4
X_17808_ net997 _02092_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_09590_ _05277_ _05279_ _05281_ _05284_ VGND VGND VPWR VPWR _05285_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08541_ CPU.rs2\[12\] _04199_ _04204_ VGND VGND VPWR VPWR _04261_ sky130_fd_sc_hd__a21o_1
X_17739_ net928 _02023_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08472_ mapped_spi_ram.div_counter\[1\] net23 _04193_ mapped_spi_ram.div_counter\[0\]
+ VGND VGND VPWR VPWR _04194_ sky130_fd_sc_hd__and4b_1
XFILLER_0_106_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_926 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09024_ _04209_ VGND VGND VPWR VPWR _04740_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_150_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15207__119 clknet_1_1__leaf__02751_ VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__inv_2
Xhold220 _01723_ VGND VGND VPWR VPWR net1461 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold231 mapped_spi_ram.state\[0\] VGND VGND VPWR VPWR net1472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 mapped_spi_flash.rcv_data\[28\] VGND VGND VPWR VPWR net1483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 mapped_spi_ram.snd_bitcount\[2\] VGND VGND VPWR VPWR net1494 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold264 mapped_spi_ram.rcv_bitcount\[0\] VGND VGND VPWR VPWR net1505 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold275 mapped_spi_ram.rbusy VGND VGND VPWR VPWR net1516 sky130_fd_sc_hd__dlygate4sd3_1
X_14924__1006 clknet_1_0__leaf__02707_ VGND VGND VPWR VPWR net1038 sky130_fd_sc_hd__inv_2
Xhold286 mapped_spi_flash.rcv_bitcount\[1\] VGND VGND VPWR VPWR net1527 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold297 CPU.state\[3\] VGND VGND VPWR VPWR net1538 sky130_fd_sc_hd__dlygate4sd3_1
X_09926_ _05552_ VGND VGND VPWR VPWR _02480_ sky130_fd_sc_hd__clkbuf_1
X_09857_ _05505_ net1853 _05491_ VGND VGND VPWR VPWR _05506_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08808_ _04524_ _04526_ _04527_ VGND VGND VPWR VPWR _04528_ sky130_fd_sc_hd__o21a_4
XTAP_TAPCELL_ROW_29_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09788_ net1812 _05008_ _05463_ VGND VGND VPWR VPWR _05465_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_104 _05401_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08739_ _04458_ _04239_ VGND VGND VPWR VPWR _04459_ sky130_fd_sc_hd__nor2_1
XANTENNA_115 _05487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_126 _05543_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_137 _05696_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_148 _07260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ mapped_spi_ram.rcv_bitcount\[0\] mapped_spi_ram.state\[3\] _06627_ VGND VGND
+ VPWR VPWR _06636_ sky130_fd_sc_hd__a21o_1
XANTENNA_159 _07302_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10701_ _06043_ VGND VGND VPWR VPWR _02149_ sky130_fd_sc_hd__clkbuf_1
X_11681_ mapped_spi_ram.rcv_data\[19\] _06588_ VGND VGND VPWR VPWR _06593_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13420_ _07841_ _07847_ _07514_ VGND VGND VPWR VPWR _07848_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_81_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14591__706 clknet_1_1__leaf__02674_ VGND VGND VPWR VPWR net738 sky130_fd_sc_hd__inv_2
X_10632_ net2399 _05996_ _06000_ _05993_ VGND VGND VPWR VPWR _02174_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_81_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13351_ CPU.registerFile\[5\]\[13\] CPU.registerFile\[4\]\[13\] net14 VGND VGND VPWR
+ VPWR _07781_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10563_ _05943_ _05957_ VGND VGND VPWR VPWR _05958_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12302_ CPU.aluIn1\[4\] _06961_ _06859_ VGND VGND VPWR VPWR _06962_ sky130_fd_sc_hd__mux2_1
X_16070_ CPU.registerFile\[15\]\[19\] CPU.registerFile\[11\]\[19\] _02849_ VGND VGND
+ VPWR VPWR _03550_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10494_ net1383 _05892_ _05902_ _05885_ VGND VGND VPWR VPWR _02214_ sky130_fd_sc_hd__o211a_1
XFILLER_0_134_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13282_ CPU.registerFile\[16\]\[11\] CPU.registerFile\[20\]\[11\] _07339_ VGND VGND
+ VPWR VPWR _07714_ sky130_fd_sc_hd__mux2_1
X_12233_ _06909_ VGND VGND VPWR VPWR _01445_ sky130_fd_sc_hd__clkbuf_1
X_15125__1155 clknet_1_1__leaf__02743_ VGND VGND VPWR VPWR net1187 sky130_fd_sc_hd__inv_2
X_12164_ CPU.aluShamt\[4\] _06854_ VGND VGND VPWR VPWR _06856_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11115_ net2240 _05691_ _06263_ VGND VGND VPWR VPWR _06264_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_112_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14411__543 clknet_1_0__leaf__02657_ VGND VGND VPWR VPWR net575 sky130_fd_sc_hd__inv_2
X_16972_ clknet_leaf_21_clk _01298_ VGND VGND VPWR VPWR CPU.mem_wdata\[3\] sky130_fd_sc_hd__dfxtp_2
X_12095_ _06818_ VGND VGND VPWR VPWR _06819_ sky130_fd_sc_hd__buf_4
X_15923_ CPU.registerFile\[5\]\[15\] CPU.registerFile\[4\]\[15\] _02806_ VGND VGND
+ VPWR VPWR _03407_ sky130_fd_sc_hd__mux2_1
X_11046_ net2507 _05691_ _06226_ VGND VGND VPWR VPWR _06227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15854_ _02771_ _03337_ _03338_ _03339_ _02807_ VGND VGND VPWR VPWR _03340_ sky130_fd_sc_hd__a221o_1
XFILLER_0_87_801 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15785_ _03268_ _03272_ _02784_ VGND VGND VPWR VPWR _03273_ sky130_fd_sc_hd__a21o_1
X_12997_ CPU.registerFile\[6\]\[3\] _07263_ VGND VGND VPWR VPWR _07437_ sky130_fd_sc_hd__or2_1
XFILLER_0_143_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17524_ net713 _01812_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_11948_ net2537 _05727_ _06733_ VGND VGND VPWR VPWR _06741_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17455_ net644 _01743_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[10\] sky130_fd_sc_hd__dfxtp_1
X_11879_ _06704_ VGND VGND VPWR VPWR _01629_ sky130_fd_sc_hd__clkbuf_1
X_16406_ _02949_ _03872_ _03875_ VGND VGND VPWR VPWR _03876_ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_119_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_156_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13618_ _08036_ _08039_ _07514_ VGND VGND VPWR VPWR _08040_ sky130_fd_sc_hd__a21oi_2
X_17386_ net575 _01674_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16337_ _02858_ _03805_ _03808_ _05029_ VGND VGND VPWR VPWR _03809_ sky130_fd_sc_hd__o211a_1
X_15076__1140 clknet_1_0__leaf__02724_ VGND VGND VPWR VPWR net1172 sky130_fd_sc_hd__inv_2
XFILLER_0_15_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13549_ CPU.registerFile\[14\]\[19\] CPU.registerFile\[10\]\[19\] _04937_ VGND VGND
+ VPWR VPWR _07973_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16268_ CPU.registerFile\[27\]\[25\] CPU.registerFile\[31\]\[25\] _02777_ VGND VGND
+ VPWR VPWR _03742_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_132_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18007_ net1180 _02287_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_15219_ clknet_1_1__leaf__02749_ VGND VGND VPWR VPWR _02753_ sky130_fd_sc_hd__buf_1
X_14039__316 clknet_1_1__leaf__08364_ VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__inv_2
X_16199_ CPU.registerFile\[22\]\[23\] _05440_ VGND VGND VPWR VPWR _03675_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14687__792 clknet_1_0__leaf__02684_ VGND VGND VPWR VPWR net824 sky130_fd_sc_hd__inv_2
X_09711_ _05401_ VGND VGND VPWR VPWR _05402_ sky130_fd_sc_hd__buf_4
X_14386__520 clknet_1_1__leaf__02655_ VGND VGND VPWR VPWR net552 sky130_fd_sc_hd__inv_2
X_09642_ _04718_ _05152_ _04636_ VGND VGND VPWR VPWR _05335_ sky130_fd_sc_hd__mux2_1
X_09573_ _05265_ _05268_ _04491_ VGND VGND VPWR VPWR _05269_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_143_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08524_ CPU.aluIn1\[21\] _04243_ VGND VGND VPWR VPWR _04244_ sky130_fd_sc_hd__or2_1
X_14085__358 clknet_1_1__leaf__08368_ VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__inv_2
XFILLER_0_78_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14852__940 clknet_1_0__leaf__02701_ VGND VGND VPWR VPWR net972 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_63_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09007_ _04476_ _04723_ VGND VGND VPWR VPWR _04724_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09909_ _05272_ VGND VGND VPWR VPWR _05541_ sky130_fd_sc_hd__buf_4
X_12920_ _07235_ VGND VGND VPWR VPWR _07361_ sky130_fd_sc_hd__buf_4
X_12851_ _07291_ _07293_ VGND VGND VPWR VPWR _07294_ sky130_fd_sc_hd__or2_1
X_11802_ _05230_ net2269 _06661_ VGND VGND VPWR VPWR _06664_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15570_ _05048_ VGND VGND VPWR VPWR _03064_ sky130_fd_sc_hd__clkbuf_4
X_11733_ mapped_spi_ram.state\[3\] _06623_ _06474_ VGND VGND VPWR VPWR _06624_ sky130_fd_sc_hd__a21o_1
XFILLER_0_139_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17240_ net430 _01528_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_11664_ net1412 _06575_ _06583_ _06581_ VGND VGND VPWR VPWR _01722_ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13403_ _07555_ _07828_ _07830_ _07831_ _07302_ VGND VGND VPWR VPWR _07832_ sky130_fd_sc_hd__a221o_1
XFILLER_0_154_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17171_ clknet_leaf_25_clk _01459_ VGND VGND VPWR VPWR CPU.mem_wmask\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10615_ net2533 _05983_ _05990_ _05980_ VGND VGND VPWR VPWR _02181_ sky130_fd_sc_hd__o211a_1
X_11595_ _06512_ _04631_ VGND VGND VPWR VPWR _06535_ sky130_fd_sc_hd__nor2_1
XFILLER_0_153_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16122_ CPU.registerFile\[12\]\[21\] _03118_ VGND VGND VPWR VPWR _03600_ sky130_fd_sc_hd__or2_1
XFILLER_0_141_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13334_ _07760_ _07761_ _07762_ _07764_ _07302_ VGND VGND VPWR VPWR _07765_ sky130_fd_sc_hd__a221o_2
XFILLER_0_134_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10546_ mapped_spi_flash.snd_bitcount\[3\] _05943_ VGND VGND VPWR VPWR _05944_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_114_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16053_ CPU.registerFile\[6\]\[19\] _02819_ VGND VGND VPWR VPWR _03533_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13265_ _07398_ _07696_ _07697_ VGND VGND VPWR VPWR _07698_ sky130_fd_sc_hd__o21a_1
Xclkbuf_1_1__f__02691_ clknet_0__02691_ VGND VGND VPWR VPWR clknet_1_1__leaf__02691_
+ sky130_fd_sc_hd__clkbuf_16
X_10477_ _04509_ _04550_ _04629_ VGND VGND VPWR VPWR _05888_ sky130_fd_sc_hd__a21oi_1
X_12216_ _06896_ VGND VGND VPWR VPWR _01449_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13196_ _07412_ _07628_ _07630_ VGND VGND VPWR VPWR _07631_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_94_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12147_ _06846_ VGND VGND VPWR VPWR _01502_ sky130_fd_sc_hd__clkbuf_1
X_16955_ net250 _01281_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_12078_ _05273_ net1855 _06805_ VGND VGND VPWR VPWR _06810_ sky130_fd_sc_hd__mux2_1
X_11029_ net1845 _05675_ _06215_ VGND VGND VPWR VPWR _06218_ sky130_fd_sc_hd__mux2_1
X_15906_ CPU.registerFile\[16\]\[14\] _02831_ _02834_ CPU.registerFile\[17\]\[14\]
+ _02854_ VGND VGND VPWR VPWR _03391_ sky130_fd_sc_hd__o221a_1
X_16886_ net2109 _04166_ _04167_ VGND VGND VPWR VPWR _02631_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15837_ CPU.registerFile\[20\]\[12\] CPU.registerFile\[21\]\[12\] _03066_ VGND VGND
+ VPWR VPWR _03324_ sky130_fd_sc_hd__mux2_1
X_15236__145 clknet_1_1__leaf__02754_ VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__inv_2
XFILLER_0_59_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15768_ CPU.registerFile\[27\]\[10\] _02928_ _02910_ VGND VGND VPWR VPWR _03257_
+ sky130_fd_sc_hd__o21a_1
X_14010__290 clknet_1_1__leaf__08361_ VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__inv_2
X_17507_ net696 _01795_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15699_ _03182_ _03189_ _02844_ VGND VGND VPWR VPWR _03190_ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14923__1005 clknet_1_0__leaf__02707_ VGND VGND VPWR VPWR net1037 sky130_fd_sc_hd__inv_2
X_17438_ net627 net1451 VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[31\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_15 _02867_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_26 _02948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_37 _03289_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_48 _04762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_133_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17369_ net558 _01657_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[1\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_59 _05007_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__08465_ clknet_0__08465_ VGND VGND VPWR VPWR clknet_1_1__leaf__08465_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_2_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_120_Left_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16649__93 clknet_1_1__leaf__03989_ VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_145_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_145_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap17 _04645_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_2
X_09625_ _04283_ _04310_ VGND VGND VPWR VPWR _05319_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_39_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09556_ _05252_ VGND VGND VPWR VPWR _05253_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_65_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15124__1154 clknet_1_0__leaf__02743_ VGND VGND VPWR VPWR net1186 sky130_fd_sc_hd__inv_2
X_08507_ CPU.rs2\[28\] _04201_ _04206_ VGND VGND VPWR VPWR _04227_ sky130_fd_sc_hd__a21o_1
XFILLER_0_148_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09487_ _04717_ _05174_ _05179_ _05186_ VGND VGND VPWR VPWR _05187_ sky130_fd_sc_hd__a211o_4
XFILLER_0_93_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_136_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10400_ _05829_ VGND VGND VPWR VPWR _02235_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11380_ _06404_ VGND VGND VPWR VPWR _01831_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14358__496 clknet_1_0__leaf__08468_ VGND VGND VPWR VPWR net528 sky130_fd_sc_hd__inv_2
XFILLER_0_150_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10331_ _05786_ VGND VGND VPWR VPWR _02262_ sky130_fd_sc_hd__clkbuf_1
X_13050_ _04971_ VGND VGND VPWR VPWR _07489_ sky130_fd_sc_hd__buf_4
X_10262_ _05749_ VGND VGND VPWR VPWR _02309_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13996__278 clknet_1_0__leaf__08359_ VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__inv_2
X_12001_ _06746_ VGND VGND VPWR VPWR _06769_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_76_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10193_ net2219 _05704_ _05692_ VGND VGND VPWR VPWR _05705_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16740_ _04050_ _04057_ _04058_ _04059_ VGND VGND VPWR VPWR _04060_ sky130_fd_sc_hd__a31o_1
X_12903_ _07252_ VGND VGND VPWR VPWR _07345_ sky130_fd_sc_hd__clkbuf_4
X_16671_ _04914_ VGND VGND VPWR VPWR _04001_ sky130_fd_sc_hd__buf_2
X_13883_ CPU.registerFile\[18\]\[30\] CPU.registerFile\[22\]\[30\] _07314_ VGND VGND
+ VPWR VPWR _08296_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14068__342 clknet_1_1__leaf__08367_ VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__inv_2
X_15622_ _02757_ _03091_ _03100_ _03114_ _02846_ VGND VGND VPWR VPWR _03115_ sky130_fd_sc_hd__a311o_2
XTAP_TAPCELL_ROW_17_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523__644 clknet_1_0__leaf__02668_ VGND VGND VPWR VPWR net676 sky130_fd_sc_hd__inv_2
X_12834_ _07238_ VGND VGND VPWR VPWR _07277_ sky130_fd_sc_hd__buf_4
XFILLER_0_33_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18341_ clknet_leaf_4_clk _02621_ VGND VGND VPWR VPWR per_uart.rx_data\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15553_ CPU.registerFile\[28\]\[5\] _02791_ VGND VGND VPWR VPWR _03047_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11716_ net1635 _06603_ _06612_ _06607_ VGND VGND VPWR VPWR _01699_ sky130_fd_sc_hd__o211a_1
X_18272_ net105 _02552_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15484_ _02813_ VGND VGND VPWR VPWR _02980_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_126_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12696_ _07177_ VGND VGND VPWR VPWR _07178_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_154_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17223_ net413 _01511_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11647_ mapped_spi_ram.rcv_bitcount\[3\] _06570_ VGND VGND VPWR VPWR _06571_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17154_ net378 _01442_ VGND VGND VPWR VPWR CPU.aluReg\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16591__62 clknet_1_0__leaf__03970_ VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__inv_2
X_11578_ net1371 _06495_ _06523_ _06516_ VGND VGND VPWR VPWR _01748_ sky130_fd_sc_hd__o211a_1
X_16105_ CPU.registerFile\[15\]\[20\] CPU.registerFile\[11\]\[20\] _02849_ VGND VGND
+ VPWR VPWR _03584_ sky130_fd_sc_hd__mux2_1
X_13317_ CPU.registerFile\[6\]\[12\] _05337_ VGND VGND VPWR VPWR _07748_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold808 CPU.registerFile\[12\]\[0\] VGND VGND VPWR VPWR net2049 sky130_fd_sc_hd__dlygate4sd3_1
X_17085_ net343 _01407_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[15\] sky130_fd_sc_hd__dfxtp_1
Xhold819 CPU.registerFile\[21\]\[13\] VGND VGND VPWR VPWR net2060 sky130_fd_sc_hd__dlygate4sd3_1
X_10529_ _05886_ _04635_ VGND VGND VPWR VPWR _05932_ sky130_fd_sc_hd__nor2_1
Xclkbuf_1_1__f__02743_ clknet_0__02743_ VGND VGND VPWR VPWR clknet_1_1__leaf__02743_
+ sky130_fd_sc_hd__clkbuf_16
X_16036_ CPU.registerFile\[6\]\[18\] _03057_ _03140_ _03516_ VGND VGND VPWR VPWR _03517_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13248_ CPU.registerFile\[18\]\[10\] CPU.registerFile\[22\]\[10\] _07315_ VGND VGND
+ VPWR VPWR _07681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__02674_ clknet_0__02674_ VGND VGND VPWR VPWR clknet_1_1__leaf__02674_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_149_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13179_ CPU.registerFile\[3\]\[8\] _04987_ _07613_ _04939_ VGND VGND VPWR VPWR _07614_
+ sky130_fd_sc_hd__o211a_1
X_17987_ clknet_leaf_7_clk net1364 VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_127_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16938_ net233 _01264_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_14606__719 clknet_1_0__leaf__02676_ VGND VGND VPWR VPWR net751 sky130_fd_sc_hd__inv_2
X_16869_ net1561 _04153_ _04155_ VGND VGND VPWR VPWR _02626_ sky130_fd_sc_hd__o21ba_1
X_09410_ _04692_ _05111_ _05112_ VGND VGND VPWR VPWR _05113_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14799__893 clknet_1_1__leaf__02695_ VGND VGND VPWR VPWR net925 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_140_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14498__621 clknet_1_0__leaf__02666_ VGND VGND VPWR VPWR net653 sky130_fd_sc_hd__inv_2
X_09341_ _05047_ VGND VGND VPWR VPWR _02568_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09272_ _04981_ VGND VGND VPWR VPWR _04982_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_118_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_603 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08987_ _04702_ _04704_ _04373_ VGND VGND VPWR VPWR _04705_ sky130_fd_sc_hd__mux2_1
Xclkbuf_2_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_3_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09608_ _04276_ _04699_ _04808_ CPU.aluReg\[6\] _05302_ VGND VGND VPWR VPWR _05303_
+ sky130_fd_sc_hd__a221o_1
X_10880_ net2056 _05731_ _06128_ VGND VGND VPWR VPWR _06138_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__02694_ clknet_0__02694_ VGND VGND VPWR VPWR clknet_1_0__leaf__02694_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09539_ _05232_ _05235_ _05112_ VGND VGND VPWR VPWR _05236_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__07221_ clknet_0__07221_ VGND VGND VPWR VPWR clknet_1_0__leaf__07221_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12550_ net1814 _05007_ _07096_ VGND VGND VPWR VPWR _07098_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11501_ CPU.mem_wmask\[1\] CPU.mem_wmask\[0\] CPU.mem_wmask\[3\] CPU.mem_wmask\[2\]
+ VGND VGND VPWR VPWR _06468_ sky130_fd_sc_hd__or4_4
X_12481_ _07061_ VGND VGND VPWR VPWR _01349_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11432_ _06431_ VGND VGND VPWR VPWR _01806_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14151_ CPU.Jimm\[19\] _08411_ _08387_ VGND VGND VPWR VPWR _08412_ sky130_fd_sc_hd__mux2_1
X_11363_ _06394_ VGND VGND VPWR VPWR _01838_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13102_ _07535_ _07538_ _07320_ VGND VGND VPWR VPWR _07539_ sky130_fd_sc_hd__mux2_2
X_10314_ _05487_ net2325 _05777_ VGND VGND VPWR VPWR _05778_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11294_ CPU.registerFile\[9\]\[0\] _05735_ _06323_ VGND VGND VPWR VPWR _06358_ sky130_fd_sc_hd__mux2_1
X_13033_ _07360_ _07468_ _07471_ _07392_ VGND VGND VPWR VPWR _07472_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_91_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17910_ net1099 net1477 VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[28\] sky130_fd_sc_hd__dfxtp_1
X_10245_ _05487_ net2155 _05740_ VGND VGND VPWR VPWR _05741_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14922__1004 clknet_1_0__leaf__02707_ VGND VGND VPWR VPWR net1036 sky130_fd_sc_hd__inv_2
X_10176_ _05693_ VGND VGND VPWR VPWR _02339_ sky130_fd_sc_hd__clkbuf_1
X_17841_ net1030 _02125_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_109_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16628__74 clknet_1_1__leaf__03971_ VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__inv_2
X_17772_ net961 _02056_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_109_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14984_ clknet_1_1__leaf__02708_ VGND VGND VPWR VPWR _02714_ sky130_fd_sc_hd__buf_1
X_16723_ _04027_ _04039_ _05175_ VGND VGND VPWR VPWR _04045_ sky130_fd_sc_hd__a21o_1
X_13935_ _07260_ _08346_ VGND VGND VPWR VPWR _08347_ sky130_fd_sc_hd__or2_1
XFILLER_0_135_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16643__88 clknet_1_1__leaf__03988_ VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__inv_2
X_13866_ _07360_ _08269_ _08272_ _08279_ VGND VGND VPWR VPWR _08280_ sky130_fd_sc_hd__a31o_1
XFILLER_0_158_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__08468_ clknet_0__08468_ VGND VGND VPWR VPWR clknet_1_0__leaf__08468_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_122_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15605_ CPU.registerFile\[25\]\[6\] _02802_ _02803_ VGND VGND VPWR VPWR _03098_ sky130_fd_sc_hd__o21a_1
X_12817_ _05337_ VGND VGND VPWR VPWR _07260_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_57_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_472 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_709 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13797_ CPU.registerFile\[19\]\[27\] _07618_ _08212_ _07417_ _07253_ VGND VGND VPWR
+ VPWR _08213_ sky130_fd_sc_hd__o221a_1
XFILLER_0_151_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15536_ CPU.registerFile\[19\]\[4\] CPU.registerFile\[17\]\[4\] _02874_ VGND VGND
+ VPWR VPWR _03031_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18324_ clknet_leaf_5_clk _02604_ VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_127_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18255_ net96 _02535_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_15467_ CPU.registerFile\[11\]\[3\] _02895_ _02911_ _02962_ VGND VGND VPWR VPWR _02963_
+ sky130_fd_sc_hd__o211a_1
X_12679_ net1502 _07166_ VGND VGND VPWR VPWR _00032_ sky130_fd_sc_hd__xor2_1
XFILLER_0_155_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17206_ net396 _01494_ VGND VGND VPWR VPWR CPU.aluShamt\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14418_ clknet_1_1__leaf__02653_ VGND VGND VPWR VPWR _02658_ sky130_fd_sc_hd__buf_1
XFILLER_0_154_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18186_ net217 _02466_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_100_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15398_ CPU.registerFile\[21\]\[1\] CPU.registerFile\[23\]\[1\] _05440_ VGND VGND
+ VPWR VPWR _02896_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17137_ net361 _01425_ VGND VGND VPWR VPWR CPU.aluReg\[1\] sky130_fd_sc_hd__dfxtp_1
Xhold605 CPU.registerFile\[13\]\[2\] VGND VGND VPWR VPWR net1846 sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 CPU.registerFile\[19\]\[25\] VGND VGND VPWR VPWR net1857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold627 CPU.registerFile\[24\]\[31\] VGND VGND VPWR VPWR net1868 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13979__262 clknet_1_1__leaf__08358_ VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__inv_2
Xhold638 CPU.registerFile\[31\]\[9\] VGND VGND VPWR VPWR net1879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold649 CPU.rs2\[20\] VGND VGND VPWR VPWR net1890 sky130_fd_sc_hd__dlygate4sd3_1
X_17068_ net326 _01390_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16019_ CPU.registerFile\[8\]\[18\] _02789_ _03117_ _03499_ VGND VGND VPWR VPWR _03500_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08910_ _04522_ _04533_ _04627_ _04629_ VGND VGND VPWR VPWR _04630_ sky130_fd_sc_hd__a31o_1
X_15123__1153 clknet_1_1__leaf__02743_ VGND VGND VPWR VPWR net1185 sky130_fd_sc_hd__inv_2
X_09890_ _05149_ VGND VGND VPWR VPWR _05528_ sky130_fd_sc_hd__buf_4
Xclkbuf_1_1__f__02657_ clknet_0__02657_ VGND VGND VPWR VPWR clknet_1_1__leaf__02657_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08841_ _04559_ _04560_ VGND VGND VPWR VPWR _04561_ sky130_fd_sc_hd__and2_1
Xclkbuf_0__02688_ _02688_ VGND VGND VPWR VPWR clknet_0__02688_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08772_ _04491_ VGND VGND VPWR VPWR _04492_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09324_ CPU.Jimm\[18\] _04812_ _04989_ CPU.cycles\[18\] VGND VGND VPWR VPWR _05031_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_157_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09255_ _04671_ _04962_ _04964_ _04678_ VGND VGND VPWR VPWR _04965_ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09186_ CPU.PC\[15\] _04844_ VGND VGND VPWR VPWR _04898_ sky130_fd_sc_hd__nand2_1
X_16570__43 clknet_1_1__leaf__03968_ VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__inv_2
XFILLER_0_31_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14552__670 clknet_1_1__leaf__02671_ VGND VGND VPWR VPWR net702 sky130_fd_sc_hd__inv_2
XFILLER_0_101_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10030_ net1802 _05027_ _05607_ VGND VGND VPWR VPWR _05610_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11981_ _04982_ net1733 _06758_ VGND VGND VPWR VPWR _06759_ sky130_fd_sc_hd__mux2_1
X_13720_ _08134_ _08135_ _08136_ _08138_ _07359_ VGND VGND VPWR VPWR _08139_ sky130_fd_sc_hd__a221o_1
X_10932_ _06166_ VGND VGND VPWR VPWR _02041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__02746_ clknet_0__02746_ VGND VGND VPWR VPWR clknet_1_0__leaf__02746_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13651_ _07351_ _08071_ VGND VGND VPWR VPWR _08072_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_104_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10863_ _06129_ VGND VGND VPWR VPWR _02073_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_27_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12602_ mapped_spi_flash.rbusy mapped_spi_ram.rbusy net1538 _05867_ VGND VGND VPWR
+ VPWR _00002_ sky130_fd_sc_hd__o31a_1
Xclkbuf_1_0__f__02677_ clknet_0__02677_ VGND VGND VPWR VPWR clknet_1_0__leaf__02677_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_27_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16370_ CPU.registerFile\[24\]\[28\] _02778_ _02780_ _03840_ VGND VGND VPWR VPWR
+ _03841_ sky130_fd_sc_hd__o211a_1
X_13582_ CPU.registerFile\[9\]\[20\] _07618_ _08004_ _07272_ _07285_ VGND VGND VPWR
+ VPWR _08005_ sky130_fd_sc_hd__o221a_1
X_10794_ _05532_ net2133 _06092_ VGND VGND VPWR VPWR _06093_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15321_ CPU.registerFile\[6\]\[0\] CPU.registerFile\[7\]\[0\] _02819_ VGND VGND VPWR
+ VPWR _02820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_137_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12533_ CPU.registerFile\[4\]\[28\] _04730_ _07085_ VGND VGND VPWR VPWR _07089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18040_ net1213 _02320_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14635__745 clknet_1_1__leaf__02679_ VGND VGND VPWR VPWR net777 sky130_fd_sc_hd__inv_2
X_15252_ clknet_1_1__leaf__02749_ VGND VGND VPWR VPWR _02756_ sky130_fd_sc_hd__buf_1
X_12464_ _07052_ VGND VGND VPWR VPWR _01357_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11415_ _05539_ net2501 _06419_ VGND VGND VPWR VPWR _06423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12395_ _04714_ net2457 _07013_ VGND VGND VPWR VPWR _07016_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14134_ _08398_ VGND VGND VPWR VPWR _01473_ sky130_fd_sc_hd__clkbuf_1
X_11346_ _05539_ net2375 _06382_ VGND VGND VPWR VPWR _06386_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14065_ clknet_1_1__leaf__08363_ VGND VGND VPWR VPWR _08367_ sky130_fd_sc_hd__buf_1
X_11277_ _06349_ VGND VGND VPWR VPWR _01879_ sky130_fd_sc_hd__clkbuf_1
X_13016_ _07230_ _07441_ _07455_ _07309_ VGND VGND VPWR VPWR _07456_ sky130_fd_sc_hd__a211o_1
X_10228_ _05728_ VGND VGND VPWR VPWR _02322_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_146_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17824_ net1013 _02108_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_10159_ net2336 _05681_ _05671_ VGND VGND VPWR VPWR _05682_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17755_ net944 _02039_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_14681__787 clknet_1_0__leaf__02683_ VGND VGND VPWR VPWR net819 sky130_fd_sc_hd__inv_2
X_14380__515 clknet_1_1__leaf__02654_ VGND VGND VPWR VPWR net547 sky130_fd_sc_hd__inv_2
X_16706_ _08457_ _04028_ _04029_ _04030_ VGND VGND VPWR VPWR _04031_ sky130_fd_sc_hd__a31o_1
X_13918_ CPU.registerFile\[5\]\[31\] _07577_ _08329_ _07638_ VGND VGND VPWR VPWR _08330_
+ sky130_fd_sc_hd__o211a_1
X_17686_ net875 _01974_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13849_ _08256_ _08263_ _04814_ VGND VGND VPWR VPWR _08264_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18307_ clknet_leaf_15_clk _02587_ VGND VGND VPWR VPWR CPU.PC\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15519_ _03012_ _03013_ _08400_ VGND VGND VPWR VPWR _03014_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09040_ _04356_ _04701_ VGND VGND VPWR VPWR _04755_ sky130_fd_sc_hd__nor2_1
X_18238_ net79 _02518_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18169_ net200 _02449_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold402 CPU.registerFile\[22\]\[15\] VGND VGND VPWR VPWR net1643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold413 CPU.registerFile\[24\]\[1\] VGND VGND VPWR VPWR net1654 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold424 CPU.registerFile\[16\]\[29\] VGND VGND VPWR VPWR net1665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 per_uart.uart0.txd_reg\[3\] VGND VGND VPWR VPWR net1676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold446 CPU.registerFile\[16\]\[23\] VGND VGND VPWR VPWR net1687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 per_uart.uart0.txd_reg\[0\] VGND VGND VPWR VPWR net1698 sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 CPU.registerFile\[2\]\[25\] VGND VGND VPWR VPWR net1709 sky130_fd_sc_hd__dlygate4sd3_1
X_09942_ _05497_ net1801 _05559_ VGND VGND VPWR VPWR _05563_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_1__f__02709_ clknet_0__02709_ VGND VGND VPWR VPWR clknet_1_1__leaf__02709_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_111_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold479 CPU.registerFile\[24\]\[4\] VGND VGND VPWR VPWR net1720 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09873_ _05516_ net1976 _05512_ VGND VGND VPWR VPWR _05517_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_5_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ CPU.aluIn1\[9\] CPU.Bimm\[9\] VGND VGND VPWR VPWR _04544_ sky130_fd_sc_hd__nor2_1
Xhold1102 CPU.registerFile\[23\]\[12\] VGND VGND VPWR VPWR net2343 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1113 CPU.registerFile\[17\]\[24\] VGND VGND VPWR VPWR net2354 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1124 CPU.registerFile\[10\]\[29\] VGND VGND VPWR VPWR net2365 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1135 CPU.registerFile\[18\]\[11\] VGND VGND VPWR VPWR net2376 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 CPU.registerFile\[27\]\[30\] VGND VGND VPWR VPWR net2387 sky130_fd_sc_hd__dlygate4sd3_1
X_08755_ _04359_ _04472_ _04474_ VGND VGND VPWR VPWR _04475_ sky130_fd_sc_hd__o21a_1
Xhold1157 CPU.registerFile\[13\]\[28\] VGND VGND VPWR VPWR net2398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1168 CPU.registerFile\[7\]\[17\] VGND VGND VPWR VPWR net2409 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1179 CPU.registerFile\[6\]\[3\] VGND VGND VPWR VPWR net2420 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_308 _07425_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08686_ _04279_ CPU.aluIn1\[5\] VGND VGND VPWR VPWR _04406_ sky130_fd_sc_hd__and2b_1
XANTENNA_319 _07914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_137_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09307_ _04339_ _04448_ VGND VGND VPWR VPWR _05015_ sky130_fd_sc_hd__xor2_2
XFILLER_0_91_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14921__1003 clknet_1_1__leaf__02707_ VGND VGND VPWR VPWR net1035 sky130_fd_sc_hd__inv_2
XFILLER_0_119_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09238_ _04242_ _04489_ _04948_ _04768_ VGND VGND VPWR VPWR _04949_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09169_ CPU.PC\[5\] CPU.Bimm\[5\] _04819_ VGND VGND VPWR VPWR _04881_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11200_ _06308_ VGND VGND VPWR VPWR _01915_ sky130_fd_sc_hd__clkbuf_1
X_12180_ _04409_ _06865_ _06868_ _06866_ _06862_ VGND VGND VPWR VPWR _01491_ sky130_fd_sc_hd__o221a_1
X_11131_ net2392 _05708_ _06263_ VGND VGND VPWR VPWR _06272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold980 CPU.registerFile\[24\]\[22\] VGND VGND VPWR VPWR net2221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold991 CPU.registerFile\[27\]\[21\] VGND VGND VPWR VPWR net2232 sky130_fd_sc_hd__dlygate4sd3_1
X_11062_ net2094 _05708_ _06226_ VGND VGND VPWR VPWR _06235_ sky130_fd_sc_hd__mux2_1
X_14216__392 clknet_1_1__leaf__08431_ VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__inv_2
X_10013_ net1774 _04748_ _05596_ VGND VGND VPWR VPWR _05601_ sky130_fd_sc_hd__mux2_1
X_15870_ _03352_ _03353_ _03355_ _02945_ VGND VGND VPWR VPWR _03356_ sky130_fd_sc_hd__o22a_2
X_16499__169 clknet_1_0__leaf__02756_ VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__inv_2
XFILLER_0_25_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17540_ net729 _01828_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_11964_ _04714_ net2284 _06747_ VGND VGND VPWR VPWR _06750_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13703_ CPU.registerFile\[16\]\[24\] CPU.registerFile\[20\]\[24\] _07648_ VGND VGND
+ VPWR VPWR _08122_ sky130_fd_sc_hd__mux2_1
X_10915_ _06157_ VGND VGND VPWR VPWR _02049_ sky130_fd_sc_hd__clkbuf_1
X_17471_ net660 _01759_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[26\] sky130_fd_sc_hd__dfxtp_1
X_11895_ _06713_ VGND VGND VPWR VPWR _01622_ sky130_fd_sc_hd__clkbuf_1
X_13634_ CPU.registerFile\[5\]\[22\] _07804_ _08054_ _07368_ VGND VGND VPWR VPWR _08055_
+ sky130_fd_sc_hd__o211a_1
X_16422_ CPU.registerFile\[26\]\[29\] _02861_ VGND VGND VPWR VPWR _03892_ sky130_fd_sc_hd__or2_1
X_10846_ _06120_ VGND VGND VPWR VPWR _02081_ sky130_fd_sc_hd__clkbuf_1
X_15122__1152 clknet_1_0__leaf__02743_ VGND VGND VPWR VPWR net1184 sky130_fd_sc_hd__inv_2
XFILLER_0_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16353_ CPU.registerFile\[25\]\[27\] _05406_ _05070_ VGND VGND VPWR VPWR _03825_
+ sky130_fd_sc_hd__o21a_1
X_13565_ CPU.registerFile\[3\]\[20\] _07804_ _07987_ VGND VGND VPWR VPWR _07988_ sky130_fd_sc_hd__o21a_1
XFILLER_0_26_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10777_ _05516_ net2248 _06081_ VGND VGND VPWR VPWR _06084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15304_ _02779_ VGND VGND VPWR VPWR _02803_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12516_ _07079_ VGND VGND VPWR VPWR _01332_ sky130_fd_sc_hd__clkbuf_1
X_16284_ CPU.registerFile\[6\]\[25\] CPU.registerFile\[7\]\[25\] _08395_ VGND VGND
+ VPWR VPWR _03758_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13496_ _07230_ _07921_ _07309_ VGND VGND VPWR VPWR _07922_ sky130_fd_sc_hd__a21o_1
X_16534__10 clknet_1_1__leaf__03965_ VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__inv_2
XFILLER_0_152_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18023_ net1196 _02303_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_12447_ _05359_ net1806 _07035_ VGND VGND VPWR VPWR _07043_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_117_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12378_ _07006_ VGND VGND VPWR VPWR _01397_ sky130_fd_sc_hd__clkbuf_1
X_14117_ _07127_ VGND VGND VPWR VPWR _08387_ sky130_fd_sc_hd__buf_4
X_11329_ _05522_ net1911 _06371_ VGND VGND VPWR VPWR _06377_ sky130_fd_sc_hd__mux2_1
X_15097_ _07187_ net1441 _02727_ VGND VGND VPWR VPWR _02278_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17807_ net996 _02091_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_15999_ CPU.registerFile\[10\]\[17\] _02816_ _02910_ VGND VGND VPWR VPWR _03481_
+ sky130_fd_sc_hd__o21a_1
X_08540_ CPU.aluIn1\[13\] _04259_ VGND VGND VPWR VPWR _04260_ sky130_fd_sc_hd__or2_1
X_17738_ net927 _02022_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_08471_ _04192_ VGND VGND VPWR VPWR _04193_ sky130_fd_sc_hd__clkbuf_4
X_17669_ net858 _01957_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14306__449 clknet_1_1__leaf__08463_ VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__inv_2
XFILLER_0_148_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09023_ _04671_ _04736_ _04738_ _04678_ VGND VGND VPWR VPWR _04739_ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_150_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold210 _01726_ VGND VGND VPWR VPWR net1451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 CPU.cycles\[6\] VGND VGND VPWR VPWR net1462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 mapped_spi_ram.rcv_data\[1\] VGND VGND VPWR VPWR net1473 sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 mapped_spi_flash.rcv_data\[17\] VGND VGND VPWR VPWR net1484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 CPU.cycles\[12\] VGND VGND VPWR VPWR net1495 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold265 mapped_spi_flash.rcv_data\[6\] VGND VGND VPWR VPWR net1506 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_53_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold276 CPU.rs2\[28\] VGND VGND VPWR VPWR net1517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 mapped_spi_flash.cmd_addr\[0\] VGND VGND VPWR VPWR net1528 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09925_ _05551_ net2181 _05533_ VGND VGND VPWR VPWR _05552_ sky130_fd_sc_hd__mux2_1
Xhold298 CPU.PC\[4\] VGND VGND VPWR VPWR net1539 sky130_fd_sc_hd__dlygate4sd3_1
X_09856_ _04797_ VGND VGND VPWR VPWR _05505_ sky130_fd_sc_hd__clkbuf_4
X_14664__771 clknet_1_1__leaf__02682_ VGND VGND VPWR VPWR net803 sky130_fd_sc_hd__inv_2
X_08807_ CPU.aluIn1\[1\] _04525_ VGND VGND VPWR VPWR _04527_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_29_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ _05464_ VGND VGND VPWR VPWR _02531_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_29_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08738_ CPU.aluIn1\[22\] VGND VGND VPWR VPWR _04458_ sky130_fd_sc_hd__inv_2
XANTENNA_105 _05401_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_116 _05487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_127 _05543_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 _05698_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08669_ CPU.aluIn1\[16\] VGND VGND VPWR VPWR _04389_ sky130_fd_sc_hd__inv_2
XANTENNA_149 _07268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_751 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10700_ _05507_ net1692 _06034_ VGND VGND VPWR VPWR _06043_ sky130_fd_sc_hd__mux2_1
X_11680_ net1610 _06590_ _06592_ _06581_ VGND VGND VPWR VPWR _01715_ sky130_fd_sc_hd__o211a_1
X_14062__337 clknet_1_1__leaf__08366_ VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__inv_2
X_10631_ mapped_spi_flash.rcv_data\[8\] _05994_ VGND VGND VPWR VPWR _06000_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_81_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13350_ _07778_ _07779_ _07476_ VGND VGND VPWR VPWR _07780_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10562_ mapped_spi_flash.snd_bitcount\[1\] mapped_spi_flash.snd_bitcount\[0\] net2543
+ VGND VGND VPWR VPWR _05957_ sky130_fd_sc_hd__o21ai_1
X_12301_ CPU.aluReg\[5\] CPU.aluReg\[3\] _06939_ VGND VGND VPWR VPWR _06961_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13281_ _07360_ _07708_ _07712_ _07380_ VGND VGND VPWR VPWR _07713_ sky130_fd_sc_hd__o211a_1
X_10493_ net1366 _05887_ _05856_ _05901_ VGND VGND VPWR VPWR _05902_ sky130_fd_sc_hd__a211o_1
X_12232_ CPU.aluReg\[21\] _06908_ _06891_ VGND VGND VPWR VPWR _06909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Left_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12163_ CPU.aluShamt\[4\] _06854_ VGND VGND VPWR VPWR _06855_ sky130_fd_sc_hd__and2_1
X_11114_ _06251_ VGND VGND VPWR VPWR _06263_ sky130_fd_sc_hd__clkbuf_4
X_14747__846 clknet_1_0__leaf__02690_ VGND VGND VPWR VPWR net878 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_112_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16971_ clknet_leaf_27_clk _01297_ VGND VGND VPWR VPWR CPU.mem_wdata\[2\] sky130_fd_sc_hd__dfxtp_2
X_12094_ _05488_ _06395_ VGND VGND VPWR VPWR _06818_ sky130_fd_sc_hd__nand2_2
X_16507__176 clknet_1_0__leaf__03962_ VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__inv_2
X_11045_ _06214_ VGND VGND VPWR VPWR _06226_ sky130_fd_sc_hd__clkbuf_4
X_15922_ _08397_ _03401_ _03405_ _02903_ VGND VGND VPWR VPWR _03406_ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15853_ CPU.registerFile\[9\]\[13\] _02778_ _03125_ VGND VGND VPWR VPWR _03339_ sky130_fd_sc_hd__o21a_1
X_15784_ _02771_ _03269_ _03270_ _03271_ _02807_ VGND VGND VPWR VPWR _03272_ sky130_fd_sc_hd__a221o_1
X_12996_ CPU.registerFile\[2\]\[3\] CPU.registerFile\[3\]\[3\] _07260_ VGND VGND VPWR
+ VPWR _07436_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Left_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17523_ net712 _01811_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11947_ _06740_ VGND VGND VPWR VPWR _01597_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17454_ net643 _01742_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11878_ CPU.registerFile\[10\]\[5\] _05725_ _06697_ VGND VGND VPWR VPWR _06704_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13617_ CPU.registerFile\[23\]\[21\] _07382_ _08038_ VGND VGND VPWR VPWR _08039_
+ sky130_fd_sc_hd__o21ai_1
X_16405_ _03227_ _03873_ _03874_ _03030_ VGND VGND VPWR VPWR _03875_ sky130_fd_sc_hd__a22o_1
X_14793__888 clknet_1_0__leaf__02694_ VGND VGND VPWR VPWR net920 sky130_fd_sc_hd__inv_2
X_10829_ _06111_ VGND VGND VPWR VPWR _02089_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_119_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17385_ net574 _01673_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14492__616 clknet_1_0__leaf__02665_ VGND VGND VPWR VPWR net648 sky130_fd_sc_hd__inv_2
XFILLER_0_144_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13548_ _07412_ _07970_ _07971_ VGND VGND VPWR VPWR _07972_ sky130_fd_sc_hd__o21a_1
X_16336_ _02818_ _03806_ _03807_ VGND VGND VPWR VPWR _03808_ sky130_fd_sc_hd__a21o_1
XFILLER_0_137_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16267_ _03739_ _03740_ _02855_ VGND VGND VPWR VPWR _03741_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13479_ _07653_ _07903_ _07904_ VGND VGND VPWR VPWR _07905_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_132_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_33_Left_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18006_ net1179 _02286_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16198_ CPU.registerFile\[21\]\[23\] CPU.registerFile\[23\]\[23\] _05440_ VGND VGND
+ VPWR VPWR _03674_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14232__407 clknet_1_0__leaf__08432_ VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__inv_2
XFILLER_0_121_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09710_ CPU.cycles\[2\] _04687_ _05388_ _05400_ VGND VGND VPWR VPWR _05401_ sky130_fd_sc_hd__a211o_2
X_14920__1002 clknet_1_1__leaf__02707_ VGND VGND VPWR VPWR net1034 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_147_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09641_ _05334_ VGND VGND VPWR VPWR _02555_ sky130_fd_sc_hd__clkbuf_1
X_09572_ _04313_ _04698_ _04218_ CPU.aluReg\[7\] _05267_ VGND VGND VPWR VPWR _05268_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08523_ CPU.rs2\[21\] _04200_ _04205_ VGND VGND VPWR VPWR _04243_ sky130_fd_sc_hd__a21o_1
XFILLER_0_148_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15213__124 clknet_1_0__leaf__02752_ VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__inv_2
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09006_ _04362_ _04467_ _04475_ VGND VGND VPWR VPWR _04723_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_689 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15121__1151 clknet_1_1__leaf__02743_ VGND VGND VPWR VPWR net1183 sky130_fd_sc_hd__inv_2
X_09908_ _05540_ VGND VGND VPWR VPWR _02486_ sky130_fd_sc_hd__clkbuf_1
X_09839_ _05493_ net1984 _05491_ VGND VGND VPWR VPWR _05494_ sky130_fd_sc_hd__mux2_1
X_12850_ CPU.registerFile\[30\]\[0\] CPU.registerFile\[26\]\[0\] _07292_ VGND VGND
+ VPWR VPWR _07293_ sky130_fd_sc_hd__mux2_1
X_11801_ _06663_ VGND VGND VPWR VPWR _01666_ sky130_fd_sc_hd__clkbuf_1
X_12781_ clknet_1_1__leaf__07223_ VGND VGND VPWR VPWR _07226_ sky130_fd_sc_hd__buf_1
XFILLER_0_69_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _06572_ _06622_ VGND VGND VPWR VPWR _06623_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15188__101 clknet_1_0__leaf__02750_ VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__inv_2
XFILLER_0_83_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14451_ clknet_1_1__leaf__02653_ VGND VGND VPWR VPWR _02661_ sky130_fd_sc_hd__buf_1
X_11663_ mapped_spi_ram.rcv_data\[27\] _06577_ VGND VGND VPWR VPWR _06583_ sky130_fd_sc_hd__or2_1
XFILLER_0_154_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_153_Right_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13402_ CPU.registerFile\[31\]\[14\] _07289_ _07290_ CPU.registerFile\[27\]\[14\]
+ _07345_ VGND VGND VPWR VPWR _07831_ sky130_fd_sc_hd__o221a_1
XFILLER_0_126_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17170_ clknet_leaf_25_clk _01458_ VGND VGND VPWR VPWR CPU.mem_wmask\[2\] sky130_fd_sc_hd__dfxtp_1
X_10614_ mapped_spi_flash.rcv_data\[15\] _05981_ VGND VGND VPWR VPWR _05990_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_12_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11594_ net1372 _06524_ _06534_ _06516_ VGND VGND VPWR VPWR _01743_ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16121_ CPU.registerFile\[14\]\[21\] CPU.registerFile\[10\]\[21\] _03082_ VGND VGND
+ VPWR VPWR _03599_ sky130_fd_sc_hd__mux2_1
X_13333_ _07351_ _07763_ VGND VGND VPWR VPWR _07764_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10545_ mapped_spi_flash.snd_bitcount\[2\] mapped_spi_flash.snd_bitcount\[1\] mapped_spi_flash.snd_bitcount\[0\]
+ VGND VGND VPWR VPWR _05943_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_114_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16052_ CPU.registerFile\[1\]\[19\] _03228_ _03531_ _02818_ VGND VGND VPWR VPWR _03532_
+ sky130_fd_sc_hd__a22o_1
X_13264_ CPU.registerFile\[13\]\[10\] _07629_ _07488_ CPU.registerFile\[9\]\[10\]
+ _07489_ VGND VGND VPWR VPWR _07697_ sky130_fd_sc_hd__o221a_1
Xclkbuf_1_1__f__02690_ clknet_0__02690_ VGND VGND VPWR VPWR clknet_1_1__leaf__02690_
+ sky130_fd_sc_hd__clkbuf_16
X_10476_ _05886_ VGND VGND VPWR VPWR _05887_ sky130_fd_sc_hd__buf_2
XFILLER_0_32_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12215_ CPU.aluReg\[25\] _06895_ _06891_ VGND VGND VPWR VPWR _06896_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13195_ CPU.registerFile\[29\]\[8\] _07629_ _07488_ CPU.registerFile\[25\]\[8\] _07489_
+ VGND VGND VPWR VPWR _07630_ sky130_fd_sc_hd__o221a_1
X_14335__475 clknet_1_1__leaf__08466_ VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_94_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12146_ _05273_ net2373 _06841_ VGND VGND VPWR VPWR _06846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13973__257 clknet_1_1__leaf__08357_ VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__inv_2
XFILLER_0_47_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16954_ net249 _01280_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_12077_ _06809_ VGND VGND VPWR VPWR _01535_ sky130_fd_sc_hd__clkbuf_1
X_11028_ _06217_ VGND VGND VPWR VPWR _01996_ sky130_fd_sc_hd__clkbuf_1
X_15905_ CPU.registerFile\[20\]\[14\] CPU.registerFile\[21\]\[14\] _03066_ VGND VGND
+ VPWR VPWR _03390_ sky130_fd_sc_hd__mux2_1
X_16885_ per_uart.uart0.rx_bitcount\[1\] per_uart.uart0.rx_bitcount\[0\] _04193_ _04137_
+ VGND VGND VPWR VPWR _04167_ sky130_fd_sc_hd__and4b_1
XFILLER_0_154_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15836_ _03319_ _03320_ _03322_ _02945_ VGND VGND VPWR VPWR _03323_ sky130_fd_sc_hd__o22a_2
XFILLER_0_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_125_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15767_ CPU.registerFile\[31\]\[10\] _03072_ VGND VGND VPWR VPWR _03256_ sky130_fd_sc_hd__or2_1
X_12979_ _07237_ VGND VGND VPWR VPWR _07420_ sky130_fd_sc_hd__buf_4
X_14801__895 clknet_1_0__leaf__02695_ VGND VGND VPWR VPWR net927 sky130_fd_sc_hd__inv_2
X_17506_ net695 _01794_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14718_ clknet_1_0__leaf__02686_ VGND VGND VPWR VPWR _02688_ sky130_fd_sc_hd__buf_1
XFILLER_0_47_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14045__321 clknet_1_1__leaf__08365_ VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__inv_2
X_15698_ _03185_ _03188_ _02809_ VGND VGND VPWR VPWR _03189_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_157_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14500__623 clknet_1_0__leaf__02666_ VGND VGND VPWR VPWR net655 sky130_fd_sc_hd__inv_2
XFILLER_0_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17437_ net626 net1408 VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[30\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_16 _02875_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_120_Right_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_27 _02948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_38 _03383_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776__225 clknet_1_1__leaf__07225_ VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__inv_2
XFILLER_0_55_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17368_ net557 _01656_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[0\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_49 _04762_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_41_Left_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16319_ CPU.registerFile\[16\]\[26\] CPU.registerFile\[18\]\[26\] _03032_ VGND VGND
+ VPWR VPWR _03792_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17299_ net488 _01587_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__08464_ clknet_0__08464_ VGND VGND VPWR VPWR clknet_1_1__leaf__08464_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_3_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_145_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_908 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09624_ _04422_ _05317_ VGND VGND VPWR VPWR _05318_ sky130_fd_sc_hd__nor2_1
Xmax_cap18 net19 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_2
XFILLER_0_69_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09555_ CPU.cycles\[8\] _04687_ _05237_ _05251_ VGND VGND VPWR VPWR _05252_ sky130_fd_sc_hd__a211o_4
XTAP_TAPCELL_ROW_65_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08506_ _04224_ _04225_ VGND VGND VPWR VPWR _04226_ sky130_fd_sc_hd__or2b_1
X_09486_ _05181_ _05185_ _04492_ VGND VGND VPWR VPWR _05186_ sky130_fd_sc_hd__o21a_1
XFILLER_0_53_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14776__872 clknet_1_0__leaf__02693_ VGND VGND VPWR VPWR net904 sky130_fd_sc_hd__inv_2
XFILLER_0_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_754 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10330_ _05507_ net2379 _05777_ VGND VGND VPWR VPWR _05786_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10261_ _05507_ net2353 _05740_ VGND VGND VPWR VPWR _05749_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12000_ _06768_ VGND VGND VPWR VPWR _01572_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_76_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10192_ _05108_ VGND VGND VPWR VPWR _05704_ sky130_fd_sc_hd__buf_2
XFILLER_0_17_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12902_ _07296_ _07343_ VGND VGND VPWR VPWR _07344_ sky130_fd_sc_hd__or2_1
X_13882_ net1523 _08018_ _08295_ _08017_ VGND VGND VPWR VPWR _01324_ sky130_fd_sc_hd__o211a_1
X_16670_ _08379_ _05375_ _08454_ VGND VGND VPWR VPWR _04000_ sky130_fd_sc_hd__or3b_1
X_14859__947 clknet_1_1__leaf__02701_ VGND VGND VPWR VPWR net979 sky130_fd_sc_hd__inv_2
X_15621_ _03106_ _03113_ _02844_ VGND VGND VPWR VPWR _03114_ sky130_fd_sc_hd__o21a_1
X_12833_ _07235_ VGND VGND VPWR VPWR _07276_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_17_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18340_ clknet_leaf_4_clk _02620_ VGND VGND VPWR VPWR per_uart.rx_data\[4\] sky130_fd_sc_hd__dfxtp_1
X_15552_ CPU.registerFile\[30\]\[5\] CPU.registerFile\[26\]\[5\] _02787_ VGND VGND
+ VPWR VPWR _03046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11715_ net1456 _06601_ VGND VGND VPWR VPWR _06612_ sky130_fd_sc_hd__or2_1
X_15483_ CPU.registerFile\[6\]\[3\] _02870_ _02894_ _02978_ VGND VGND VPWR VPWR _02979_
+ sky130_fd_sc_hd__o211a_1
X_18271_ net104 _02551_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_12695_ per_uart.tx_busy per_uart.uart0.tx_wr VGND VGND VPWR VPWR _07177_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_154_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17222_ net412 _01510_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11646_ mapped_spi_ram.rcv_bitcount\[2\] mapped_spi_ram.rcv_bitcount\[1\] mapped_spi_ram.rcv_bitcount\[0\]
+ VGND VGND VPWR VPWR _06570_ sky130_fd_sc_hd__or3_1
XFILLER_0_80_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17153_ net377 _01441_ VGND VGND VPWR VPWR CPU.aluReg\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11577_ net1386 _06517_ _06509_ _06522_ VGND VGND VPWR VPWR _06523_ sky130_fd_sc_hd__a211o_1
XFILLER_0_123_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13316_ CPU.registerFile\[2\]\[12\] CPU.registerFile\[3\]\[12\] _07260_ VGND VGND
+ VPWR VPWR _07747_ sky130_fd_sc_hd__mux2_1
X_16104_ _03195_ _03580_ _03581_ _03582_ _03245_ VGND VGND VPWR VPWR _03583_ sky130_fd_sc_hd__a221o_1
X_17084_ net342 _01406_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_10528_ net1354 _05892_ _05931_ _05885_ VGND VGND VPWR VPWR _02209_ sky130_fd_sc_hd__o211a_1
X_14296_ clknet_1_0__leaf__08433_ VGND VGND VPWR VPWR _08463_ sky130_fd_sc_hd__buf_1
Xhold809 CPU.registerFile\[24\]\[11\] VGND VGND VPWR VPWR net2050 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13247_ _07254_ _07675_ _07679_ _07646_ VGND VGND VPWR VPWR _07680_ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16035_ CPU.registerFile\[7\]\[18\] _03317_ VGND VGND VPWR VPWR _03516_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10459_ _05852_ _05872_ VGND VGND VPWR VPWR _05873_ sky130_fd_sc_hd__nor2_1
Xclkbuf_1_1__f__02673_ clknet_0__02673_ VGND VGND VPWR VPWR clknet_1_1__leaf__02673_
+ sky130_fd_sc_hd__clkbuf_16
X_15242__150 clknet_1_1__leaf__02755_ VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__inv_2
X_13178_ CPU.registerFile\[2\]\[8\] _07388_ VGND VGND VPWR VPWR _07613_ sky130_fd_sc_hd__or2_1
X_12129_ _05109_ net1836 _06830_ VGND VGND VPWR VPWR _06837_ sky130_fd_sc_hd__mux2_1
X_17986_ net1174 _02270_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_16937_ net232 _01263_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_127_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16868_ per_uart.uart0.rx_count16\[0\] per_uart.uart0.rx_busy _08355_ _04589_ VGND
+ VGND VPWR VPWR _04155_ sky130_fd_sc_hd__a31o_1
X_15819_ _02771_ _03303_ _03304_ _03305_ _02807_ VGND VGND VPWR VPWR _03306_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_36_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16799_ _04803_ _04914_ _03990_ VGND VGND VPWR VPWR _04109_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_140_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_140_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09340_ CPU.registerFile\[16\]\[18\] _05046_ _04983_ VGND VGND VPWR VPWR _05047_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09271_ _04969_ _04973_ _04980_ VGND VGND VPWR VPWR _04981_ sky130_fd_sc_hd__or3b_4
XFILLER_0_74_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15120__1150 clknet_1_1__leaf__02743_ VGND VGND VPWR VPWR net1182 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_60_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f__03989_ clknet_0__03989_ VGND VGND VPWR VPWR clknet_1_1__leaf__03989_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_99_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15040__1109 clknet_1_0__leaf__02718_ VGND VGND VPWR VPWR net1141 sky130_fd_sc_hd__inv_2
X_13956__241 clknet_1_0__leaf__08356_ VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__inv_2
XFILLER_0_139_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08986_ _04477_ _04703_ VGND VGND VPWR VPWR _04704_ sky130_fd_sc_hd__and2b_1
X_14017__297 clknet_1_0__leaf__08361_ VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__inv_2
XFILLER_0_3_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14210__387 clknet_1_1__leaf__08430_ VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_3_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09607_ CPU.aluIn1\[6\] _04274_ _04698_ VGND VGND VPWR VPWR _05302_ sky130_fd_sc_hd__and3_1
Xclkbuf_1_0__f__02693_ clknet_0__02693_ VGND VGND VPWR VPWR clknet_1_0__leaf__02693_
+ sky130_fd_sc_hd__clkbuf_16
X_09538_ _05234_ VGND VGND VPWR VPWR _05235_ sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__07220_ clknet_0__07220_ VGND VGND VPWR VPWR clknet_1_0__leaf__07220_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_94_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09469_ _05169_ VGND VGND VPWR VPWR _05170_ sky130_fd_sc_hd__buf_4
XFILLER_0_149_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11500_ _06467_ VGND VGND VPWR VPWR _01774_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12480_ net1796 _05691_ _07060_ VGND VGND VPWR VPWR _07061_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11431_ _05555_ net2196 _06396_ VGND VGND VPWR VPWR _06431_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14150_ _08410_ VGND VGND VPWR VPWR _08411_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_78_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11362_ _05555_ net1876 _06359_ VGND VGND VPWR VPWR _06394_ sky130_fd_sc_hd__mux2_1
X_13101_ CPU.registerFile\[21\]\[6\] _07244_ _07429_ CPU.registerFile\[17\]\[6\] _07537_
+ VGND VGND VPWR VPWR _07538_ sky130_fd_sc_hd__o221a_1
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10313_ _05776_ VGND VGND VPWR VPWR _05777_ sky130_fd_sc_hd__buf_4
XFILLER_0_104_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11293_ _06357_ VGND VGND VPWR VPWR _01871_ sky130_fd_sc_hd__clkbuf_1
X_13032_ CPU.registerFile\[1\]\[4\] _07387_ _07470_ _07231_ VGND VGND VPWR VPWR _07471_
+ sky130_fd_sc_hd__a211o_1
X_10244_ _05739_ VGND VGND VPWR VPWR _05740_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_91_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17840_ net1029 _02124_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_10175_ net2154 _05691_ _05692_ VGND VGND VPWR VPWR _05693_ sky130_fd_sc_hd__mux2_1
X_17771_ net960 _02055_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_109_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16722_ _03991_ net1820 VGND VGND VPWR VPWR _04044_ sky130_fd_sc_hd__nand2_1
X_13934_ CPU.registerFile\[28\]\[31\] CPU.registerFile\[24\]\[31\] _04936_ VGND VGND
+ VPWR VPWR _08346_ sky130_fd_sc_hd__mux2_1
X_14447__576 clknet_1_0__leaf__02660_ VGND VGND VPWR VPWR net608 sky130_fd_sc_hd__inv_2
XFILLER_0_135_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13865_ _08275_ _08278_ _07474_ VGND VGND VPWR VPWR _08279_ sky130_fd_sc_hd__a21oi_2
X_14185__364 clknet_1_1__leaf__08428_ VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__08467_ clknet_0__08467_ VGND VGND VPWR VPWR clknet_1_0__leaf__08467_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_122_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15604_ CPU.registerFile\[29\]\[6\] _02800_ VGND VGND VPWR VPWR _03097_ sky130_fd_sc_hd__or2_1
X_12816_ CPU.registerFile\[1\]\[0\] _07256_ _07257_ _07258_ VGND VGND VPWR VPWR _07259_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_922 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13796_ CPU.registerFile\[18\]\[27\] CPU.registerFile\[22\]\[27\] _07457_ VGND VGND
+ VPWR VPWR _08212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18323_ clknet_leaf_15_clk _02603_ VGND VGND VPWR VPWR CPU.PC\[23\] sky130_fd_sc_hd__dfxtp_1
X_15535_ _02939_ VGND VGND VPWR VPWR _03030_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_151_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18254_ net95 _02534_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15466_ CPU.registerFile\[15\]\[3\] _02826_ VGND VGND VPWR VPWR _02962_ sky130_fd_sc_hd__or2_1
X_12678_ _07166_ _07167_ VGND VGND VPWR VPWR _00031_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17205_ net395 net1543 VGND VGND VPWR VPWR CPU.aluShamt\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11629_ _06551_ _06557_ _06499_ VGND VGND VPWR VPWR _06558_ sky130_fd_sc_hd__o21ai_1
X_18185_ net216 _02465_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_100_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15397_ _02894_ VGND VGND VPWR VPWR _02895_ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_7_Left_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_874 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14913__996 clknet_1_0__leaf__02706_ VGND VGND VPWR VPWR net1028 sky130_fd_sc_hd__inv_2
XFILLER_0_52_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17136_ net360 _01424_ VGND VGND VPWR VPWR CPU.aluReg\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold606 CPU.registerFile\[2\]\[15\] VGND VGND VPWR VPWR net1847 sky130_fd_sc_hd__dlygate4sd3_1
Xhold617 CPU.registerFile\[7\]\[1\] VGND VGND VPWR VPWR net1858 sky130_fd_sc_hd__dlygate4sd3_1
X_14612__724 clknet_1_0__leaf__02677_ VGND VGND VPWR VPWR net756 sky130_fd_sc_hd__inv_2
Xhold628 CPU.registerFile\[20\]\[16\] VGND VGND VPWR VPWR net1869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold639 CPU.registerFile\[14\]\[11\] VGND VGND VPWR VPWR net1880 sky130_fd_sc_hd__dlygate4sd3_1
X_14279_ _08457_ _05418_ VGND VGND VPWR VPWR _08458_ sky130_fd_sc_hd__nor2_1
X_17067_ net325 _01389_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16018_ CPU.registerFile\[12\]\[18\] _03118_ VGND VGND VPWR VPWR _03499_ sky130_fd_sc_hd__or2_1
Xclkbuf_0__02756_ _02756_ VGND VGND VPWR VPWR clknet_0__02756_ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f__02656_ clknet_0__02656_ VGND VGND VPWR VPWR clknet_1_1__leaf__02656_
+ sky130_fd_sc_hd__clkbuf_16
X_08840_ CPU.aluIn1\[16\] _04494_ VGND VGND VPWR VPWR _04560_ sky130_fd_sc_hd__or2_1
Xclkbuf_0__02687_ _02687_ VGND VGND VPWR VPWR clknet_0__02687_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08771_ CPU.instr\[2\] _04196_ VGND VGND VPWR VPWR _04491_ sky130_fd_sc_hd__nor2_2
X_17969_ net1157 _02253_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_0_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09323_ _04782_ _05029_ _04777_ VGND VGND VPWR VPWR _05030_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_149_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_903 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09254_ _04670_ _04963_ VGND VGND VPWR VPWR _04964_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09185_ CPU.PC\[14\] _04846_ _04896_ VGND VGND VPWR VPWR _04897_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_141_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14888__973 clknet_1_1__leaf__02704_ VGND VGND VPWR VPWR net1005 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_73_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08969_ net19 VGND VGND VPWR VPWR _04688_ sky130_fd_sc_hd__buf_4
X_11980_ _06746_ VGND VGND VPWR VPWR _06758_ sky130_fd_sc_hd__buf_4
X_10931_ net1604 _05712_ _06165_ VGND VGND VPWR VPWR _06166_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__02745_ clknet_0__02745_ VGND VGND VPWR VPWR clknet_1_0__leaf__02745_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_98_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10862_ net2176 _05712_ _06128_ VGND VGND VPWR VPWR _06129_ sky130_fd_sc_hd__mux2_1
X_13650_ CPU.registerFile\[30\]\[22\] CPU.registerFile\[26\]\[22\] _07297_ VGND VGND
+ VPWR VPWR _08071_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_104_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__02676_ clknet_0__02676_ VGND VGND VPWR VPWR clknet_1_0__leaf__02676_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_27_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12601_ _05813_ _06014_ _06030_ VGND VGND VPWR VPWR _00005_ sky130_fd_sc_hd__a21oi_1
X_13581_ CPU.registerFile\[8\]\[20\] CPU.registerFile\[12\]\[20\] _07339_ VGND VGND
+ VPWR VPWR _08004_ sky130_fd_sc_hd__mux2_1
X_10793_ _06069_ VGND VGND VPWR VPWR _06092_ sky130_fd_sc_hd__clkbuf_4
X_12532_ _07088_ VGND VGND VPWR VPWR _01292_ sky130_fd_sc_hd__clkbuf_1
X_15320_ _08394_ VGND VGND VPWR VPWR _02819_ sky130_fd_sc_hd__buf_4
XFILLER_0_94_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12463_ net2075 _05675_ _07049_ VGND VGND VPWR VPWR _07052_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14202_ clknet_1_0__leaf__08363_ VGND VGND VPWR VPWR _08430_ sky130_fd_sc_hd__buf_1
X_11414_ _06422_ VGND VGND VPWR VPWR _01815_ sky130_fd_sc_hd__clkbuf_1
X_12394_ _07015_ VGND VGND VPWR VPWR _01390_ sky130_fd_sc_hd__clkbuf_1
X_14133_ CPU.Jimm\[15\] _08397_ _08387_ VGND VGND VPWR VPWR _08398_ sky130_fd_sc_hd__mux2_1
X_11345_ _06385_ VGND VGND VPWR VPWR _01847_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11276_ CPU.registerFile\[9\]\[9\] _05717_ _06346_ VGND VGND VPWR VPWR _06349_ sky130_fd_sc_hd__mux2_1
X_13015_ _07271_ _07444_ _07447_ _07454_ _07306_ VGND VGND VPWR VPWR _07455_ sky130_fd_sc_hd__o311a_1
X_10227_ net2281 _05727_ _05713_ VGND VGND VPWR VPWR _05728_ sky130_fd_sc_hd__mux2_1
X_17823_ net1012 _02107_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_10158_ _04761_ VGND VGND VPWR VPWR _05681_ sky130_fd_sc_hd__buf_2
XFILLER_0_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17754_ net943 _02038_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_10089_ _05641_ VGND VGND VPWR VPWR _02374_ sky130_fd_sc_hd__clkbuf_1
X_16705_ _03995_ _05245_ _07123_ VGND VGND VPWR VPWR _04030_ sky130_fd_sc_hd__o21ai_1
X_13917_ CPU.registerFile\[4\]\[31\] _07291_ VGND VGND VPWR VPWR _08329_ sky130_fd_sc_hd__or2_1
X_17685_ net874 _01973_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13848_ _07379_ _08258_ _08262_ _07268_ VGND VGND VPWR VPWR _08263_ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13779_ _07474_ _08192_ _08195_ VGND VGND VPWR VPWR _08196_ sky130_fd_sc_hd__or3_1
XFILLER_0_57_465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18306_ clknet_leaf_15_clk _02586_ VGND VGND VPWR VPWR CPU.PC\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15518_ CPU.registerFile\[30\]\[4\] CPU.registerFile\[26\]\[4\] _02881_ VGND VGND
+ VPWR VPWR _03013_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_702 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18237_ net78 _02517_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_15449_ _02938_ _02941_ _02944_ _02945_ VGND VGND VPWR VPWR _02946_ sky130_fd_sc_hd__o22a_1
XFILLER_0_53_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18168_ net199 _02448_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_135_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold403 CPU.registerFile\[10\]\[26\] VGND VGND VPWR VPWR net1644 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold414 CPU.registerFile\[30\]\[18\] VGND VGND VPWR VPWR net1655 sky130_fd_sc_hd__dlygate4sd3_1
X_17119_ clknet_leaf_18_clk _00021_ VGND VGND VPWR VPWR CPU.cycles\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold425 CPU.registerFile\[20\]\[22\] VGND VGND VPWR VPWR net1666 sky130_fd_sc_hd__dlygate4sd3_1
X_18099_ net162 _02379_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[29\] sky130_fd_sc_hd__dfxtp_1
Xhold436 CPU.registerFile\[16\]\[17\] VGND VGND VPWR VPWR net1677 sky130_fd_sc_hd__dlygate4sd3_1
Xhold447 CPU.registerFile\[4\]\[24\] VGND VGND VPWR VPWR net1688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 CPU.registerFile\[14\]\[30\] VGND VGND VPWR VPWR net1699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 CPU.registerFile\[5\]\[22\] VGND VGND VPWR VPWR net1710 sky130_fd_sc_hd__dlygate4sd3_1
X_09941_ _05562_ VGND VGND VPWR VPWR _02475_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_1__f__02708_ clknet_0__02708_ VGND VGND VPWR VPWR clknet_1_1__leaf__02708_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_55_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ _05026_ VGND VGND VPWR VPWR _05516_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_5_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ _04542_ _04516_ _04515_ _04513_ VGND VGND VPWR VPWR _04543_ sky130_fd_sc_hd__a31oi_4
Xhold1103 CPU.registerFile\[21\]\[28\] VGND VGND VPWR VPWR net2344 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1114 CPU.registerFile\[19\]\[15\] VGND VGND VPWR VPWR net2355 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1125 CPU.registerFile\[11\]\[31\] VGND VGND VPWR VPWR net2366 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1136 CPU.registerFile\[20\]\[25\] VGND VGND VPWR VPWR net2377 sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ _04473_ _04229_ VGND VGND VPWR VPWR _04474_ sky130_fd_sc_hd__or2_1
Xhold1147 CPU.registerFile\[6\]\[6\] VGND VGND VPWR VPWR net2388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1158 mapped_spi_flash.rcv_data\[7\] VGND VGND VPWR VPWR net2399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 CPU.registerFile\[27\]\[1\] VGND VGND VPWR VPWR net2410 sky130_fd_sc_hd__dlygate4sd3_1
X_14983__1059 clknet_1_1__leaf__02713_ VGND VGND VPWR VPWR net1091 sky130_fd_sc_hd__inv_2
X_08685_ _04274_ CPU.aluIn1\[6\] VGND VGND VPWR VPWR _04405_ sky130_fd_sc_hd__and2b_1
XANTENNA_309 _07653_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09306_ _04449_ _05013_ VGND VGND VPWR VPWR _05014_ sky130_fd_sc_hd__and2_1
XFILLER_0_137_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09237_ _04945_ _04947_ _04374_ VGND VGND VPWR VPWR _04948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_134_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09168_ _04867_ _04869_ _04878_ _04879_ VGND VGND VPWR VPWR _04880_ sky130_fd_sc_hd__a31o_1
XFILLER_0_133_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09099_ _04805_ _04807_ _04810_ _04491_ VGND VGND VPWR VPWR _04811_ sky130_fd_sc_hd__o31a_1
XFILLER_0_102_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11130_ _06271_ VGND VGND VPWR VPWR _01948_ sky130_fd_sc_hd__clkbuf_1
Xhold970 CPU.registerFile\[26\]\[29\] VGND VGND VPWR VPWR net2211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 per_uart.uart0.tx_wr VGND VGND VPWR VPWR net2222 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_79_Left_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11061_ _06234_ VGND VGND VPWR VPWR _01980_ sky130_fd_sc_hd__clkbuf_1
Xhold992 CPU.registerFile\[25\]\[22\] VGND VGND VPWR VPWR net2233 sky130_fd_sc_hd__dlygate4sd3_1
X_10012_ _05600_ VGND VGND VPWR VPWR _02410_ sky130_fd_sc_hd__clkbuf_1
X_14751_ clknet_1_1__leaf__02686_ VGND VGND VPWR VPWR _02691_ sky130_fd_sc_hd__buf_1
XFILLER_0_25_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11963_ _06749_ VGND VGND VPWR VPWR _01590_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14641__750 clknet_1_0__leaf__02680_ VGND VGND VPWR VPWR net782 sky130_fd_sc_hd__inv_2
XFILLER_0_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_86_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ _07273_ _08119_ _08120_ VGND VGND VPWR VPWR _08121_ sky130_fd_sc_hd__o21ai_2
X_10914_ net1701 _05696_ _06154_ VGND VGND VPWR VPWR _06157_ sky130_fd_sc_hd__mux2_1
X_17470_ net659 _01758_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[25\] sky130_fd_sc_hd__dfxtp_1
X_11894_ net1669 _05673_ _06711_ VGND VGND VPWR VPWR _06713_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_88_Left_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16421_ CPU.registerFile\[28\]\[29\] CPU.registerFile\[24\]\[29\] _02761_ VGND VGND
+ VPWR VPWR _03891_ sky130_fd_sc_hd__mux2_1
X_13633_ CPU.registerFile\[4\]\[22\] _07374_ VGND VGND VPWR VPWR _08054_ sky130_fd_sc_hd__or2_1
X_10845_ net2370 _05696_ _06117_ VGND VGND VPWR VPWR _06120_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__02659_ clknet_0__02659_ VGND VGND VPWR VPWR clknet_1_0__leaf__02659_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16352_ CPU.registerFile\[29\]\[27\] _03064_ VGND VGND VPWR VPWR _03824_ sky130_fd_sc_hd__or2_1
X_13564_ _04938_ VGND VGND VPWR VPWR _07987_ sky130_fd_sc_hd__clkbuf_4
X_10776_ _06083_ VGND VGND VPWR VPWR _02114_ sky130_fd_sc_hd__clkbuf_1
X_14559__677 clknet_1_0__leaf__02671_ VGND VGND VPWR VPWR net709 sky130_fd_sc_hd__inv_2
XFILLER_0_137_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15303_ _02777_ VGND VGND VPWR VPWR _02802_ sky130_fd_sc_hd__buf_4
X_12515_ net2125 _05727_ _07071_ VGND VGND VPWR VPWR _07079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16283_ CPU.registerFile\[1\]\[25\] _02873_ _03756_ _08404_ VGND VGND VPWR VPWR _03757_
+ sky130_fd_sc_hd__a22o_1
X_13495_ _07914_ _07920_ _07514_ VGND VGND VPWR VPWR _07921_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18022_ net1195 _02302_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_12446_ _07042_ VGND VGND VPWR VPWR _01365_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_676 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12377_ _05333_ net2162 _06999_ VGND VGND VPWR VPWR _07006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14116_ _08386_ VGND VGND VPWR VPWR _01467_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_97_Left_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11328_ _06376_ VGND VGND VPWR VPWR _01855_ sky130_fd_sc_hd__clkbuf_1
X_15096_ per_uart.uart0.enable16_counter\[7\] _07185_ net1440 VGND VGND VPWR VPWR
+ _02735_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_157_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11259_ CPU.registerFile\[9\]\[17\] _05700_ _06335_ VGND VGND VPWR VPWR _06340_ sky130_fd_sc_hd__mux2_1
X_14724__825 clknet_1_1__leaf__02688_ VGND VGND VPWR VPWR net857 sky130_fd_sc_hd__inv_2
X_17806_ net995 _02090_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_15998_ CPU.registerFile\[14\]\[17\] _02889_ VGND VGND VPWR VPWR _03480_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_50_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17737_ net926 _02021_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08470_ net2 VGND VGND VPWR VPWR _04192_ sky130_fd_sc_hd__clkbuf_4
X_17668_ net857 _01956_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16619_ net1797 net1591 _03979_ VGND VGND VPWR VPWR _03985_ sky130_fd_sc_hd__mux2_1
X_17599_ net788 _01887_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09022_ _04360_ _04737_ _04671_ VGND VGND VPWR VPWR _04738_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_14_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14770__867 clknet_1_1__leaf__02692_ VGND VGND VPWR VPWR net899 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_150_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold200 _02735_ VGND VGND VPWR VPWR net1441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16530__197 clknet_1_0__leaf__03964_ VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__inv_2
XFILLER_0_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold211 mapped_spi_flash.snd_bitcount\[3\] VGND VGND VPWR VPWR net1452 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_890 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold222 mapped_spi_ram.rcv_data\[28\] VGND VGND VPWR VPWR net1463 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold233 mapped_spi_ram.snd_bitcount\[4\] VGND VGND VPWR VPWR net1474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 CPU.cycles\[19\] VGND VGND VPWR VPWR net1485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 CPU.cycles\[8\] VGND VGND VPWR VPWR net1496 sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 mapped_spi_flash.snd_bitcount\[1\] VGND VGND VPWR VPWR net1507 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 mapped_spi_ram.rcv_bitcount\[4\] VGND VGND VPWR VPWR net1518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 per_uart.uart0.tx_count16\[0\] VGND VGND VPWR VPWR net1529 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09924_ _05401_ VGND VGND VPWR VPWR _05551_ sky130_fd_sc_hd__buf_4
Xhold299 per_uart.uart0.rxd_reg\[1\] VGND VGND VPWR VPWR net1540 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09855_ _05504_ VGND VGND VPWR VPWR _02503_ sky130_fd_sc_hd__clkbuf_1
X_08806_ CPU.aluIn1\[1\] _04525_ VGND VGND VPWR VPWR _04526_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_147_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09786_ net2229 _04982_ _05463_ VGND VGND VPWR VPWR _05464_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14363__500 clknet_1_0__leaf__02652_ VGND VGND VPWR VPWR net532 sky130_fd_sc_hd__inv_2
X_14939__1019 clknet_1_0__leaf__02709_ VGND VGND VPWR VPWR net1051 sky130_fd_sc_hd__inv_2
X_08737_ _04452_ _04456_ _04242_ VGND VGND VPWR VPWR _04457_ sky130_fd_sc_hd__a21oi_2
XPHY_EDGE_ROW_134_Right_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_106 _05402_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_117 _05487_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_128 _05543_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08668_ CPU.aluIn1\[17\] _04251_ VGND VGND VPWR VPWR _04388_ sky130_fd_sc_hd__and2_1
XANTENNA_139 _05698_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_101_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08599_ _04318_ _04269_ _04267_ _04264_ VGND VGND VPWR VPWR _04319_ sky130_fd_sc_hd__a31o_1
XFILLER_0_49_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10630_ net2505 _05996_ _05999_ _05993_ VGND VGND VPWR VPWR _02175_ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10561_ net1452 _05950_ _05952_ _05956_ VGND VGND VPWR VPWR _02201_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12300_ _06960_ VGND VGND VPWR VPWR _01429_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13280_ _07369_ _07709_ _07711_ _07231_ VGND VGND VPWR VPWR _07712_ sky130_fd_sc_hd__a211o_1
XFILLER_0_51_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10492_ _05886_ _05900_ VGND VGND VPWR VPWR _05901_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12231_ CPU.aluIn1\[21\] _06907_ _06894_ VGND VGND VPWR VPWR _06908_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12162_ CPU.aluShamt\[3\] CPU.aluShamt\[2\] CPU.aluShamt\[1\] CPU.aluShamt\[0\] VGND
+ VGND VPWR VPWR _06854_ sky130_fd_sc_hd__or4_1
XFILLER_0_20_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11113_ _06262_ VGND VGND VPWR VPWR _01956_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16970_ clknet_leaf_22_clk _01296_ VGND VGND VPWR VPWR CPU.mem_wdata\[1\] sky130_fd_sc_hd__dfxtp_2
X_12093_ _06817_ VGND VGND VPWR VPWR _01527_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_112_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11044_ _06225_ VGND VGND VPWR VPWR _01988_ sky130_fd_sc_hd__clkbuf_1
X_15921_ _03195_ _03402_ _03404_ _02965_ VGND VGND VPWR VPWR _03405_ sky130_fd_sc_hd__a211o_1
X_15852_ CPU.registerFile\[13\]\[13\] _03123_ VGND VGND VPWR VPWR _03338_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15783_ CPU.registerFile\[9\]\[11\] _02778_ _03125_ VGND VGND VPWR VPWR _03271_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12995_ CPU.registerFile\[1\]\[3\] _07256_ _07434_ _07258_ VGND VGND VPWR VPWR _07435_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17522_ net711 _01810_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_11946_ CPU.registerFile\[11\]\[5\] _05725_ _06733_ VGND VGND VPWR VPWR _06740_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16598__69 clknet_1_1__leaf__03970_ VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__inv_2
X_17453_ net642 _01741_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[8\] sky130_fd_sc_hd__dfxtp_1
X_11877_ _06703_ VGND VGND VPWR VPWR _01630_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16404_ CPU.registerFile\[19\]\[29\] CPU.registerFile\[17\]\[29\] _03025_ VGND VGND
+ VPWR VPWR _03874_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13616_ CPU.registerFile\[19\]\[21\] _07503_ _08037_ _07296_ _07278_ VGND VGND VPWR
+ VPWR _08038_ sky130_fd_sc_hd__o221a_1
X_17384_ net573 _01672_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_10828_ net1787 _05679_ _06106_ VGND VGND VPWR VPWR _06111_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_119_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14596_ clknet_1_1__leaf__02675_ VGND VGND VPWR VPWR _02676_ sky130_fd_sc_hd__buf_1
XFILLER_0_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16335_ CPU.registerFile\[2\]\[27\] _02821_ _02822_ CPU.registerFile\[3\]\[27\] _02874_
+ VGND VGND VPWR VPWR _03807_ sky130_fd_sc_hd__a221o_1
X_13547_ CPU.registerFile\[13\]\[19\] _07414_ _07326_ CPU.registerFile\[9\]\[19\]
+ _07489_ VGND VGND VPWR VPWR _07971_ sky130_fd_sc_hd__o221a_1
XFILLER_0_55_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10759_ _06074_ VGND VGND VPWR VPWR _02122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16266_ CPU.registerFile\[28\]\[25\] CPU.registerFile\[24\]\[25\] _02772_ VGND VGND
+ VPWR VPWR _03740_ sky130_fd_sc_hd__mux2_1
X_13478_ CPU.registerFile\[13\]\[17\] _07281_ _07404_ CPU.registerFile\[9\]\[17\]
+ _04972_ VGND VGND VPWR VPWR _07904_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_132_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14982__1058 clknet_1_1__leaf__02713_ VGND VGND VPWR VPWR net1090 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_132_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18005_ net1178 _00007_ VGND VGND VPWR VPWR mapped_spi_flash.state\[3\] sky130_fd_sc_hd__dfxtp_1
X_12429_ _07033_ VGND VGND VPWR VPWR _01373_ sky130_fd_sc_hd__clkbuf_1
X_16197_ CPU.registerFile\[19\]\[23\] CPU.registerFile\[17\]\[23\] _02874_ VGND VGND
+ VPWR VPWR _03673_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15079_ net1363 net1341 VGND VGND VPWR VPWR _02725_ sky130_fd_sc_hd__nand2_1
X_14312__454 clknet_1_1__leaf__08464_ VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_147_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09640_ net1886 _05333_ _05189_ VGND VGND VPWR VPWR _05334_ sky130_fd_sc_hd__mux2_1
X_13950__236 clknet_1_0__leaf__07226_ VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__inv_2
X_09571_ _04210_ _05266_ _04273_ VGND VGND VPWR VPWR _05267_ sky130_fd_sc_hd__o21a_1
X_08522_ _04240_ _04241_ VGND VGND VPWR VPWR _04242_ sky130_fd_sc_hd__nor2_2
XFILLER_0_78_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09005_ _04228_ _04214_ _04681_ CPU.aluReg\[28\] _04721_ VGND VGND VPWR VPWR _04722_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09907_ _05539_ net2401 _05533_ VGND VGND VPWR VPWR _05540_ sky130_fd_sc_hd__mux2_1
X_14287__431 clknet_1_0__leaf__08462_ VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__inv_2
X_09838_ _04695_ VGND VGND VPWR VPWR _05493_ sky130_fd_sc_hd__clkbuf_4
X_09769_ net1735 _04714_ _05452_ VGND VGND VPWR VPWR _05455_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11800_ _05209_ net2036 _06661_ VGND VGND VPWR VPWR _06663_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_83_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11731_ mapped_spi_ram.rcv_bitcount\[4\] _06571_ mapped_spi_ram.rcv_bitcount\[5\]
+ VGND VGND VPWR VPWR _06622_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11662_ net1460 _06575_ _06582_ _06581_ VGND VGND VPWR VPWR _01723_ sky130_fd_sc_hd__o211a_1
X_13401_ _07296_ _07829_ VGND VGND VPWR VPWR _07830_ sky130_fd_sc_hd__or2_1
X_10613_ net2330 _05983_ _05989_ _05980_ VGND VGND VPWR VPWR _02182_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_12_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11593_ net1359 _06517_ _06509_ _06533_ VGND VGND VPWR VPWR _06534_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_12_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14753__851 clknet_1_0__leaf__02691_ VGND VGND VPWR VPWR net883 sky130_fd_sc_hd__inv_2
XFILLER_0_52_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16120_ CPU.aluIn1\[20\] _02958_ _03579_ _03598_ _02995_ VGND VGND VPWR VPWR _02434_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_24_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13332_ CPU.registerFile\[28\]\[12\] CPU.registerFile\[24\]\[12\] _07352_ VGND VGND
+ VPWR VPWR _07763_ sky130_fd_sc_hd__mux2_1
X_10544_ _05825_ _05941_ _05942_ VGND VGND VPWR VPWR _02204_ sky130_fd_sc_hd__o21a_1
X_16513__181 clknet_1_0__leaf__03963_ VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__inv_2
XFILLER_0_134_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16051_ CPU.registerFile\[5\]\[19\] CPU.registerFile\[4\]\[19\] _05092_ VGND VGND
+ VPWR VPWR _03531_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13263_ CPU.registerFile\[8\]\[10\] CPU.registerFile\[12\]\[10\] _07265_ VGND VGND
+ VPWR VPWR _07696_ sky130_fd_sc_hd__mux2_1
X_10475_ _05817_ VGND VGND VPWR VPWR _05886_ sky130_fd_sc_hd__buf_2
XFILLER_0_134_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12214_ CPU.aluIn1\[25\] _06893_ _06894_ VGND VGND VPWR VPWR _06895_ sky130_fd_sc_hd__mux2_1
X_13194_ _07234_ VGND VGND VPWR VPWR _07629_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_94_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12145_ _06845_ VGND VGND VPWR VPWR _01503_ sky130_fd_sc_hd__clkbuf_1
X_16953_ net248 _01279_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_12076_ _05253_ net1926 _06805_ VGND VGND VPWR VPWR _06809_ sky130_fd_sc_hd__mux2_1
X_15904_ _03385_ _03386_ _03388_ _02945_ VGND VGND VPWR VPWR _03389_ sky130_fd_sc_hd__o22a_2
X_11027_ net2015 _05673_ _06215_ VGND VGND VPWR VPWR _06217_ sky130_fd_sc_hd__mux2_1
X_16884_ per_uart.uart0.rx_bitcount\[0\] _04164_ _04166_ VGND VGND VPWR VPWR _02630_
+ sky130_fd_sc_hd__o21a_1
X_17480__26 VGND VGND VPWR VPWR _17480__26/HI net26 sky130_fd_sc_hd__conb_1
XFILLER_0_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15835_ CPU.registerFile\[1\]\[12\] _02939_ _03321_ _02943_ VGND VGND VPWR VPWR _03322_
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_29_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15766_ CPU.registerFile\[25\]\[10\] CPU.registerFile\[29\]\[10\] _03254_ VGND VGND
+ VPWR VPWR _03255_ sky130_fd_sc_hd__mux2_1
X_12978_ CPU.registerFile\[8\]\[2\] CPU.registerFile\[12\]\[2\] _07315_ VGND VGND
+ VPWR VPWR _07419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17505_ net694 _01793_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_142_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11929_ CPU.registerFile\[11\]\[13\] _05708_ _06722_ VGND VGND VPWR VPWR _06731_
+ sky130_fd_sc_hd__mux2_1
X_15697_ _02827_ _03186_ _03187_ VGND VGND VPWR VPWR _03188_ sky130_fd_sc_hd__o21ai_1
X_14836__926 clknet_1_0__leaf__02699_ VGND VGND VPWR VPWR net958 sky130_fd_sc_hd__inv_2
XFILLER_0_86_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17436_ net625 _01724_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_17 _02887_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_28 _02956_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17367_ net556 _01655_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[31\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_39 _03530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16318_ CPU.registerFile\[19\]\[26\] CPU.registerFile\[17\]\[26\] _02874_ VGND VGND
+ VPWR VPWR _03791_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_86 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17298_ net487 _01586_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__08463_ clknet_0__08463_ VGND VGND VPWR VPWR clknet_1_1__leaf__08463_
+ sky130_fd_sc_hd__clkbuf_16
X_14938__1018 clknet_1_0__leaf__02709_ VGND VGND VPWR VPWR net1050 sky130_fd_sc_hd__inv_2
X_16249_ _02775_ _03722_ _03723_ VGND VGND VPWR VPWR _03724_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14882__968 clknet_1_1__leaf__02703_ VGND VGND VPWR VPWR net1000 sky130_fd_sc_hd__inv_2
XFILLER_0_128_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09623_ _04282_ _04420_ _04421_ VGND VGND VPWR VPWR _05317_ sky130_fd_sc_hd__nor3_1
Xmax_cap19 _04614_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_39_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09554_ _04974_ _05239_ _05241_ _04955_ _05250_ VGND VGND VPWR VPWR _05251_ sky130_fd_sc_hd__o221ai_4
XTAP_TAPCELL_ROW_65_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08505_ CPU.aluIn1\[29\] _04223_ VGND VGND VPWR VPWR _04225_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09485_ _04323_ _04489_ _05184_ _04679_ VGND VGND VPWR VPWR _05185_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14475__601 clknet_1_1__leaf__02663_ VGND VGND VPWR VPWR net633 sky130_fd_sc_hd__inv_2
XFILLER_0_136_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10260_ _05748_ VGND VGND VPWR VPWR _02310_ sky130_fd_sc_hd__clkbuf_1
X_10191_ _05703_ VGND VGND VPWR VPWR _02334_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_76_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12901_ CPU.registerFile\[30\]\[1\] CPU.registerFile\[26\]\[1\] _07297_ VGND VGND
+ VPWR VPWR _07343_ sky130_fd_sc_hd__mux2_1
X_13881_ _07394_ _08280_ _08294_ _08015_ VGND VGND VPWR VPWR _08295_ sky130_fd_sc_hd__a211o_1
X_15620_ _03109_ _03112_ _02809_ VGND VGND VPWR VPWR _03113_ sky130_fd_sc_hd__a21oi_4
X_12832_ CPU.registerFile\[14\]\[0\] CPU.registerFile\[10\]\[0\] _07274_ VGND VGND
+ VPWR VPWR _07275_ sky130_fd_sc_hd__mux2_1
X_14981__1057 clknet_1_1__leaf__02713_ VGND VGND VPWR VPWR net1089 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _03040_ _03044_ _02784_ VGND VGND VPWR VPWR _03045_ sky130_fd_sc_hd__a21o_1
XFILLER_0_139_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11714_ net1456 _06603_ _06611_ _06607_ VGND VGND VPWR VPWR _01700_ sky130_fd_sc_hd__o211a_1
X_18270_ net103 _02550_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_15482_ CPU.registerFile\[7\]\[3\] _05092_ VGND VGND VPWR VPWR _02978_ sky130_fd_sc_hd__or2_1
X_12694_ net1426 _07174_ VGND VGND VPWR VPWR _00039_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17221_ net411 _01509_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_14341__480 clknet_1_0__leaf__08467_ VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__inv_2
X_11645_ net1332 mapped_spi_ram.state\[3\] VGND VGND VPWR VPWR _06569_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17152_ net376 _01440_ VGND VGND VPWR VPWR CPU.aluReg\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11576_ _06512_ _05906_ VGND VGND VPWR VPWR _06522_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16103_ CPU.registerFile\[10\]\[20\] _02928_ _02910_ VGND VGND VPWR VPWR _03582_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_96_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13315_ CPU.registerFile\[1\]\[12\] _07256_ _07745_ _07258_ VGND VGND VPWR VPWR _07746_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17083_ net341 _01405_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_10527_ net1402 _05887_ _05856_ _05930_ VGND VGND VPWR VPWR _05931_ sky130_fd_sc_hd__a211o_1
X_16034_ _03510_ _03514_ _03138_ VGND VGND VPWR VPWR _03515_ sky130_fd_sc_hd__a21o_1
X_13246_ _07639_ _07676_ _07677_ _07678_ _07570_ VGND VGND VPWR VPWR _07679_ sky130_fd_sc_hd__a221o_1
X_10458_ CPU.PC\[15\] _05867_ _05870_ _05871_ VGND VGND VPWR VPWR _05872_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_0_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__02672_ clknet_0__02672_ VGND VGND VPWR VPWR clknet_1_1__leaf__02672_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_149_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13177_ CPU.registerFile\[6\]\[8\] CPU.registerFile\[7\]\[8\] _07371_ VGND VGND VPWR
+ VPWR _07612_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10389_ mapped_spi_flash.snd_bitcount\[4\] mapped_spi_flash.snd_bitcount\[3\] mapped_spi_flash.snd_bitcount\[2\]
+ _05818_ VGND VGND VPWR VPWR _05819_ sky130_fd_sc_hd__or4_1
X_12128_ _06836_ VGND VGND VPWR VPWR _01511_ sky130_fd_sc_hd__clkbuf_1
X_17985_ net1173 _02269_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_12059_ _05090_ net1779 _06794_ VGND VGND VPWR VPWR _06800_ sky130_fd_sc_hd__mux2_1
X_16936_ clknet_leaf_7_clk _01262_ VGND VGND VPWR VPWR per_uart.uart0.txd_reg\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_127_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16867_ net1515 _06482_ _07195_ _04154_ VGND VGND VPWR VPWR _02625_ sky130_fd_sc_hd__a31o_1
X_12782__230 clknet_1_1__leaf__07226_ VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__inv_2
X_15818_ CPU.registerFile\[9\]\[12\] _02778_ _03125_ VGND VGND VPWR VPWR _03305_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16798_ _04052_ _04930_ _08453_ VGND VGND VPWR VPWR _04108_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_36_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_140_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14424__555 clknet_1_0__leaf__02658_ VGND VGND VPWR VPWR net587 sky130_fd_sc_hd__inv_2
X_15749_ CPU.registerFile\[19\]\[10\] CPU.registerFile\[17\]\[10\] _03025_ VGND VGND
+ VPWR VPWR _03238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09270_ _04974_ _04975_ _04978_ _04955_ _04979_ VGND VGND VPWR VPWR _04980_ sky130_fd_sc_hd__o221a_1
XFILLER_0_8_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17419_ net608 _01707_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_60_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__03988_ clknet_0__03988_ VGND VGND VPWR VPWR clknet_1_1__leaf__03988_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_155_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_9_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14470__597 clknet_1_1__leaf__02662_ VGND VGND VPWR VPWR net629 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_58_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08985_ _04226_ _04380_ _04476_ VGND VGND VPWR VPWR _04703_ sky130_fd_sc_hd__or3_1
XFILLER_0_139_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09606_ _04277_ _04806_ VGND VGND VPWR VPWR _05301_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14245__418 clknet_1_1__leaf__08434_ VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__02692_ clknet_0__02692_ VGND VGND VPWR VPWR clknet_1_0__leaf__02692_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09537_ mapped_spi_ram.rcv_data\[16\] _04645_ _05233_ VGND VGND VPWR VPWR _05234_
+ sky130_fd_sc_hd__a21oi_1
X_14819__910 clknet_1_0__leaf__02698_ VGND VGND VPWR VPWR net942 sky130_fd_sc_hd__inv_2
XFILLER_0_149_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14399__532 clknet_1_0__leaf__02656_ VGND VGND VPWR VPWR net564 sky130_fd_sc_hd__inv_2
X_09468_ _05154_ _05156_ _05168_ VGND VGND VPWR VPWR _05169_ sky130_fd_sc_hd__or3_4
XFILLER_0_19_530 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09399_ _04672_ _05100_ _05102_ _04679_ VGND VGND VPWR VPWR _05103_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11430_ _06430_ VGND VGND VPWR VPWR _01807_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_22_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11361_ _06393_ VGND VGND VPWR VPWR _01839_ sky130_fd_sc_hd__clkbuf_1
X_10312_ _05775_ _05738_ VGND VGND VPWR VPWR _05776_ sky130_fd_sc_hd__nand2_4
X_13100_ _07245_ _07536_ VGND VGND VPWR VPWR _07537_ sky130_fd_sc_hd__or2_1
X_11292_ CPU.registerFile\[9\]\[1\] _05733_ _06323_ VGND VGND VPWR VPWR _06357_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Left_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13031_ CPU.registerFile\[5\]\[4\] _04987_ _07469_ _07368_ VGND VGND VPWR VPWR _07470_
+ sky130_fd_sc_hd__o211a_1
X_10243_ _05737_ _05738_ VGND VGND VPWR VPWR _05739_ sky130_fd_sc_hd__nand2_4
XFILLER_0_30_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14865__952 clknet_1_0__leaf__02702_ VGND VGND VPWR VPWR net984 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_91_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10174_ _05670_ VGND VGND VPWR VPWR _05692_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17770_ net959 _02054_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_109_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16721_ _04038_ _04043_ _04015_ VGND VGND VPWR VPWR _02590_ sky130_fd_sc_hd__a21oi_1
X_13933_ _07519_ _08343_ _08344_ VGND VGND VPWR VPWR _08345_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13864_ _07650_ _08276_ _08277_ VGND VGND VPWR VPWR _08278_ sky130_fd_sc_hd__o21ai_1
X_14937__1017 clknet_1_0__leaf__02709_ VGND VGND VPWR VPWR net1049 sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__08466_ clknet_0__08466_ VGND VGND VPWR VPWR clknet_1_0__leaf__08466_
+ sky130_fd_sc_hd__clkbuf_16
X_15603_ CPU.registerFile\[27\]\[6\] CPU.registerFile\[31\]\[6\] _03050_ VGND VGND
+ VPWR VPWR _03096_ sky130_fd_sc_hd__mux2_1
X_12815_ _05284_ VGND VGND VPWR VPWR _07258_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_122_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13795_ CPU.registerFile\[1\]\[27\] _07387_ _08210_ _07379_ VGND VGND VPWR VPWR _08211_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_97_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18322_ clknet_leaf_15_clk _02602_ VGND VGND VPWR VPWR CPU.PC\[22\] sky130_fd_sc_hd__dfxtp_2
X_15534_ _03022_ _03023_ _03024_ _03027_ _03028_ VGND VGND VPWR VPWR _03029_ sky130_fd_sc_hd__o221a_1
X_12746_ clknet_1_0__leaf__07220_ VGND VGND VPWR VPWR _07221_ sky130_fd_sc_hd__buf_1
XFILLER_0_57_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_606 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18253_ net94 _02533_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_15465_ _02959_ _02960_ _02875_ VGND VGND VPWR VPWR _02961_ sky130_fd_sc_hd__mux2_1
X_12677_ net1447 _07164_ VGND VGND VPWR VPWR _07167_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17204_ net394 _01492_ VGND VGND VPWR VPWR CPU.aluShamt\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18184_ net215 _02464_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_11628_ mapped_spi_ram.snd_bitcount\[4\] _06550_ VGND VGND VPWR VPWR _06557_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15396_ _05406_ VGND VGND VPWR VPWR _02894_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_100_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17135_ clknet_leaf_25_clk net1427 VGND VGND VPWR VPWR CPU.cycles\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11559_ _06508_ VGND VGND VPWR VPWR _06509_ sky130_fd_sc_hd__buf_2
Xhold607 CPU.registerFile\[29\]\[18\] VGND VGND VPWR VPWR net1848 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold618 CPU.registerFile\[30\]\[4\] VGND VGND VPWR VPWR net1859 sky130_fd_sc_hd__dlygate4sd3_1
X_17066_ net324 _01388_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[28\] sky130_fd_sc_hd__dfxtp_1
Xhold629 CPU.registerFile\[17\]\[26\] VGND VGND VPWR VPWR net1870 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__02724_ clknet_0__02724_ VGND VGND VPWR VPWR clknet_1_1__leaf__02724_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14278_ _05289_ VGND VGND VPWR VPWR _08457_ sky130_fd_sc_hd__buf_2
XFILLER_0_150_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16017_ CPU.registerFile\[14\]\[18\] CPU.registerFile\[10\]\[18\] _03082_ VGND VGND
+ VPWR VPWR _03498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_761 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13229_ CPU.registerFile\[31\]\[9\] _07482_ _07420_ CPU.registerFile\[27\]\[9\] _07483_
+ VGND VGND VPWR VPWR _07663_ sky130_fd_sc_hd__o221a_1
Xclkbuf_0__02755_ _02755_ VGND VGND VPWR VPWR clknet_0__02755_ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f__02655_ clknet_0__02655_ VGND VGND VPWR VPWR clknet_1_1__leaf__02655_
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_0__02686_ _02686_ VGND VGND VPWR VPWR clknet_0__02686_ sky130_fd_sc_hd__clkbuf_16
X_08770_ _04376_ _04486_ _04489_ _04370_ VGND VGND VPWR VPWR _04490_ sky130_fd_sc_hd__a2bb2o_1
X_17968_ net1156 _02252_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_16919_ CPU.mem_wdata\[5\] _04180_ _04188_ _04176_ VGND VGND VPWR VPWR _02643_ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17899_ net1088 net1455 VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[17\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_108_Left_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09322_ mapped_spi_ram.rcv_data\[10\] _04783_ _04784_ mapped_spi_flash.rcv_data\[10\]
+ VGND VGND VPWR VPWR _05029_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_158_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_157_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09253_ _04345_ _04451_ VGND VGND VPWR VPWR _04963_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09184_ CPU.PC\[14\] _04846_ _04895_ VGND VGND VPWR VPWR _04896_ sky130_fd_sc_hd__a21o_1
X_15249__157 clknet_1_0__leaf__02755_ VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__inv_2
XFILLER_0_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_117_Left_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14980__1056 clknet_1_1__leaf__02713_ VGND VGND VPWR VPWR net1088 sky130_fd_sc_hd__inv_2
X_14587__702 clknet_1_0__leaf__02674_ VGND VGND VPWR VPWR net734 sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__08429_ clknet_0__08429_ VGND VGND VPWR VPWR clknet_1_1__leaf__08429_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_73_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08968_ _04502_ VGND VGND VPWR VPWR _04687_ sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_126_Left_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08899_ mapped_spi_ram.rcv_data\[7\] net19 _04618_ mapped_spi_flash.rcv_data\[7\]
+ VGND VGND VPWR VPWR _04619_ sky130_fd_sc_hd__a22oi_4
X_10930_ _06142_ VGND VGND VPWR VPWR _06165_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_0__f__02744_ clknet_0__02744_ VGND VGND VPWR VPWR clknet_1_0__leaf__02744_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10861_ _06105_ VGND VGND VPWR VPWR _06128_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_104_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__02675_ clknet_0__02675_ VGND VGND VPWR VPWR clknet_1_0__leaf__02675_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12600_ net1472 _06471_ _05942_ VGND VGND VPWR VPWR _00010_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_27_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13580_ _07818_ _08001_ _08002_ VGND VGND VPWR VPWR _08003_ sky130_fd_sc_hd__o21a_1
XFILLER_0_109_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10792_ _06091_ VGND VGND VPWR VPWR _02106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12531_ net1572 _04713_ _07085_ VGND VGND VPWR VPWR _07088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_135_Left_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12462_ _07051_ VGND VGND VPWR VPWR _01358_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11413_ _05537_ net2468 _06419_ VGND VGND VPWR VPWR _06422_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12393_ _04696_ net2016 _07013_ VGND VGND VPWR VPWR _07015_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14132_ _08396_ VGND VGND VPWR VPWR _08397_ sky130_fd_sc_hd__buf_4
XFILLER_0_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11344_ _05537_ CPU.registerFile\[23\]\[9\] _06382_ VGND VGND VPWR VPWR _06385_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14453__581 clknet_1_0__leaf__02661_ VGND VGND VPWR VPWR net613 sky130_fd_sc_hd__inv_2
XFILLER_0_39_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11275_ _06348_ VGND VGND VPWR VPWR _01880_ sky130_fd_sc_hd__clkbuf_1
X_13014_ _07288_ _07450_ _07452_ _07453_ _07302_ VGND VGND VPWR VPWR _07454_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_148_Right_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10226_ _05358_ VGND VGND VPWR VPWR _05727_ sky130_fd_sc_hd__clkbuf_4
X_10157_ _05680_ VGND VGND VPWR VPWR _02345_ sky130_fd_sc_hd__clkbuf_1
X_17822_ net1011 _02106_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_17753_ net942 _02037_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_10088_ net2397 _04798_ _05633_ VGND VGND VPWR VPWR _05641_ sky130_fd_sc_hd__mux2_1
X_13916_ _07801_ _08325_ _08326_ _08327_ _07555_ VGND VGND VPWR VPWR _08328_ sky130_fd_sc_hd__a221o_1
X_16704_ _08379_ _05241_ _04006_ VGND VGND VPWR VPWR _04029_ sky130_fd_sc_hd__or3b_1
X_17684_ net873 _01972_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_13847_ _07638_ _08259_ _08260_ _08261_ _07554_ VGND VGND VPWR VPWR _08262_ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16566_ clknet_1_1__leaf__07219_ VGND VGND VPWR VPWR _03968_ sky130_fd_sc_hd__buf_1
XFILLER_0_71_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13778_ _07418_ _08193_ _08194_ VGND VGND VPWR VPWR _08195_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18305_ clknet_leaf_13_clk _02585_ VGND VGND VPWR VPWR CPU.PC\[5\] sky130_fd_sc_hd__dfxtp_1
X_15517_ CPU.registerFile\[28\]\[4\] CPU.registerFile\[24\]\[4\] _02881_ VGND VGND
+ VPWR VPWR _03012_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12729_ per_uart.d_in_uart\[4\] _07178_ _07203_ per_uart.uart0.txd_reg\[5\] VGND
+ VGND VPWR VPWR _07209_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_139_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18236_ net77 _02516_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15448_ _02758_ VGND VGND VPWR VPWR _02945_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18167_ net198 _02447_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_14536__656 clknet_1_0__leaf__02669_ VGND VGND VPWR VPWR net688 sky130_fd_sc_hd__inv_2
XFILLER_0_111_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15379_ _08405_ _02871_ _02876_ VGND VGND VPWR VPWR _02877_ sky130_fd_sc_hd__a21o_1
XFILLER_0_111_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17118_ clknet_leaf_18_clk _00020_ VGND VGND VPWR VPWR CPU.cycles\[14\] sky130_fd_sc_hd__dfxtp_1
Xhold404 CPU.registerFile\[22\]\[26\] VGND VGND VPWR VPWR net1645 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold415 CPU.mem_wdata\[0\] VGND VGND VPWR VPWR net1656 sky130_fd_sc_hd__dlygate4sd3_1
X_18098_ net161 _02378_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[28\] sky130_fd_sc_hd__dfxtp_1
Xhold426 CPU.registerFile\[5\]\[29\] VGND VGND VPWR VPWR net1667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 CPU.registerFile\[28\]\[1\] VGND VGND VPWR VPWR net1678 sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 CPU.registerFile\[12\]\[14\] VGND VGND VPWR VPWR net1689 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold459 CPU.registerFile\[5\]\[31\] VGND VGND VPWR VPWR net1700 sky130_fd_sc_hd__dlygate4sd3_1
X_09940_ _05495_ net1690 _05559_ VGND VGND VPWR VPWR _05562_ sky130_fd_sc_hd__mux2_1
X_17049_ net307 _01371_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[11\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__02707_ clknet_0__02707_ VGND VGND VPWR VPWR clknet_1_1__leaf__02707_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_111_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_115_Right_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09871_ _05515_ VGND VGND VPWR VPWR _02498_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ CPU.aluIn1\[7\] CPU.Bimm\[7\] _04538_ _04541_ _04539_ VGND VGND VPWR VPWR
+ _04542_ sky130_fd_sc_hd__a221o_1
Xclkbuf_0__02669_ _02669_ VGND VGND VPWR VPWR clknet_0__02669_ sky130_fd_sc_hd__clkbuf_16
Xhold1104 CPU.registerFile\[23\]\[25\] VGND VGND VPWR VPWR net2345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1115 CPU.registerFile\[2\]\[13\] VGND VGND VPWR VPWR net2356 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1126 CPU.registerFile\[10\]\[8\] VGND VGND VPWR VPWR net2367 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 mapped_spi_ram.rcv_data\[7\] VGND VGND VPWR VPWR net2378 sky130_fd_sc_hd__dlygate4sd3_1
X_08753_ CPU.aluIn1\[27\] VGND VGND VPWR VPWR _04473_ sky130_fd_sc_hd__inv_2
Xhold1148 CPU.registerFile\[21\]\[0\] VGND VGND VPWR VPWR net2389 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 CPU.registerFile\[27\]\[29\] VGND VGND VPWR VPWR net2400 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14582__698 clknet_1_1__leaf__02673_ VGND VGND VPWR VPWR net730 sky130_fd_sc_hd__inv_2
X_08684_ _04272_ CPU.aluIn1\[7\] VGND VGND VPWR VPWR _04404_ sky130_fd_sc_hd__and2b_1
XFILLER_0_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09305_ _04448_ _04387_ _04446_ VGND VGND VPWR VPWR _05013_ sky130_fd_sc_hd__or3_1
XFILLER_0_63_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09236_ _04457_ _04946_ VGND VGND VPWR VPWR _04947_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09167_ CPU.PC\[4\] _04866_ VGND VGND VPWR VPWR _04879_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09098_ _04348_ _04699_ _04808_ CPU.aluReg\[23\] _04809_ VGND VGND VPWR VPWR _04810_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14936__1016 clknet_1_0__leaf__02709_ VGND VGND VPWR VPWR net1048 sky130_fd_sc_hd__inv_2
Xhold960 CPU.registerFile\[26\]\[17\] VGND VGND VPWR VPWR net2201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 CPU.registerFile\[17\]\[5\] VGND VGND VPWR VPWR net2212 sky130_fd_sc_hd__dlygate4sd3_1
X_11060_ net2116 _05706_ _06226_ VGND VGND VPWR VPWR _06234_ sky130_fd_sc_hd__mux2_1
Xhold982 CPU.registerFile\[14\]\[4\] VGND VGND VPWR VPWR net2223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold993 CPU.registerFile\[1\]\[8\] VGND VGND VPWR VPWR net2234 sky130_fd_sc_hd__dlygate4sd3_1
X_10011_ net1907 _04731_ _05596_ VGND VGND VPWR VPWR _05600_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11962_ _04696_ net1932 _06747_ VGND VGND VPWR VPWR _06749_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13701_ CPU.registerFile\[23\]\[24\] _07361_ _07283_ CPU.registerFile\[19\]\[24\]
+ _07253_ VGND VGND VPWR VPWR _08120_ sky130_fd_sc_hd__o221a_1
X_10913_ _06156_ VGND VGND VPWR VPWR _02050_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_86_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11893_ _06712_ VGND VGND VPWR VPWR _01623_ sky130_fd_sc_hd__clkbuf_1
X_16420_ _03015_ _03887_ _03888_ _03889_ _02930_ VGND VGND VPWR VPWR _03890_ sky130_fd_sc_hd__a221o_1
X_13632_ _07801_ _08050_ _08051_ _08052_ _07555_ VGND VGND VPWR VPWR _08053_ sky130_fd_sc_hd__a221o_1
XFILLER_0_156_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10844_ _06119_ VGND VGND VPWR VPWR _02082_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_143_Left_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__02658_ clknet_0__02658_ VGND VGND VPWR VPWR clknet_1_0__leaf__02658_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16351_ CPU.registerFile\[27\]\[27\] CPU.registerFile\[31\]\[27\] _02851_ VGND VGND
+ VPWR VPWR _03823_ sky130_fd_sc_hd__mux2_1
X_13563_ CPU.registerFile\[2\]\[20\] _07322_ VGND VGND VPWR VPWR _07986_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10775_ _05514_ net1980 _06081_ VGND VGND VPWR VPWR _06083_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15302_ CPU.registerFile\[29\]\[0\] _02800_ VGND VGND VPWR VPWR _02801_ sky130_fd_sc_hd__or2_1
X_12514_ _07078_ VGND VGND VPWR VPWR _01333_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16282_ CPU.registerFile\[5\]\[25\] CPU.registerFile\[4\]\[25\] _02805_ VGND VGND
+ VPWR VPWR _03756_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_907 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13494_ _07917_ _07919_ _07320_ VGND VGND VPWR VPWR _07920_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18021_ net1194 _02301_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12445_ _05333_ net1922 _07035_ VGND VGND VPWR VPWR _07042_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_117_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12376_ _07005_ VGND VGND VPWR VPWR _01398_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14115_ _04664_ _05212_ _00000_ VGND VGND VPWR VPWR _08386_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11327_ _05520_ net2426 _06371_ VGND VGND VPWR VPWR _06376_ sky130_fd_sc_hd__mux2_1
X_15095_ _07186_ _02734_ _02727_ VGND VGND VPWR VPWR _02277_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_152_Left_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11258_ _06339_ VGND VGND VPWR VPWR _01888_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10209_ net2003 _05715_ _05713_ VGND VGND VPWR VPWR _05716_ sky130_fd_sc_hd__mux2_1
X_11189_ _05518_ net2326 _06299_ VGND VGND VPWR VPWR _06303_ sky130_fd_sc_hd__mux2_1
X_17805_ net994 _02089_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_15997_ CPU.registerFile\[8\]\[17\] CPU.registerFile\[12\]\[17\] _02999_ VGND VGND
+ VPWR VPWR _03479_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17736_ net925 _02020_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17667_ net856 _01955_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16618_ _03984_ VGND VGND VPWR VPWR _02546_ sky130_fd_sc_hd__clkbuf_1
X_17598_ net787 _01886_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[16\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09021_ _04359_ _04232_ _04357_ VGND VGND VPWR VPWR _04737_ sky130_fd_sc_hd__nor3_1
X_18219_ net60 _02499_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold201 mapped_spi_flash.cmd_addr\[2\] VGND VGND VPWR VPWR net1442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 mapped_spi_flash.rcv_data\[29\] VGND VGND VPWR VPWR net1453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 per_uart.uart0.enable16_counter\[5\] VGND VGND VPWR VPWR net1464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 mapped_spi_flash.rcv_data\[24\] VGND VGND VPWR VPWR net1475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 mapped_spi_flash.rcv_data\[4\] VGND VGND VPWR VPWR net1486 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold256 _07145_ VGND VGND VPWR VPWR net1497 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold267 per_uart.uart0.rxd_reg\[0\] VGND VGND VPWR VPWR net1508 sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 per_uart.uart0.rx_ack VGND VGND VPWR VPWR net1519 sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ _05550_ VGND VGND VPWR VPWR _02481_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold289 CPU.rs2\[22\] VGND VGND VPWR VPWR net1530 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09854_ _05503_ net1759 _05491_ VGND VGND VPWR VPWR _05504_ sky130_fd_sc_hd__mux2_1
X_08805_ CPU.Iimm\[1\] CPU.Bimm\[1\] CPU.instr\[5\] VGND VGND VPWR VPWR _04525_ sky130_fd_sc_hd__mux2_4
X_09785_ _05451_ VGND VGND VPWR VPWR _05463_ sky130_fd_sc_hd__buf_4
XFILLER_0_147_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14699__803 clknet_1_1__leaf__02685_ VGND VGND VPWR VPWR net835 sky130_fd_sc_hd__inv_2
X_08736_ _04453_ _04243_ _04455_ VGND VGND VPWR VPWR _04456_ sky130_fd_sc_hd__o21ba_1
XANTENNA_107 _05402_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_118 _05511_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_129 _05545_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08667_ _04386_ _04249_ VGND VGND VPWR VPWR _04387_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_68_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08598_ _04314_ _04273_ _04271_ _04316_ _04317_ VGND VGND VPWR VPWR _04318_ sky130_fd_sc_hd__a311o_1
XFILLER_0_95_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_81_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10560_ _05944_ _05955_ VGND VGND VPWR VPWR _05956_ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14519__640 clknet_1_1__leaf__02668_ VGND VGND VPWR VPWR net672 sky130_fd_sc_hd__inv_2
XFILLER_0_51_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09219_ _04818_ _04913_ _04916_ _04930_ VGND VGND VPWR VPWR _04931_ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18371__30 VGND VGND VPWR VPWR _18371__30/HI net30 sky130_fd_sc_hd__conb_1
XFILLER_0_106_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10491_ CPU.PC\[10\] _05867_ _05899_ net1285 VGND VGND VPWR VPWR _05900_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_133_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12230_ CPU.aluReg\[22\] CPU.aluReg\[20\] _06906_ VGND VGND VPWR VPWR _06907_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12161_ _06853_ VGND VGND VPWR VPWR _01495_ sky130_fd_sc_hd__clkbuf_1
X_11112_ net2264 _05689_ _06252_ VGND VGND VPWR VPWR _06262_ sky130_fd_sc_hd__mux2_1
X_12092_ _05448_ net1742 _06782_ VGND VGND VPWR VPWR _06817_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_112_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold790 CPU.registerFile\[7\]\[18\] VGND VGND VPWR VPWR net2031 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11043_ net1668 _05689_ _06215_ VGND VGND VPWR VPWR _06225_ sky130_fd_sc_hd__mux2_1
X_15920_ CPU.registerFile\[15\]\[15\] _02826_ _02770_ _03403_ VGND VGND VPWR VPWR
+ _03404_ sky130_fd_sc_hd__o211a_1
X_15851_ CPU.registerFile\[15\]\[13\] CPU.registerFile\[11\]\[13\] _02906_ VGND VGND
+ VPWR VPWR _03337_ sky130_fd_sc_hd__mux2_1
X_14565__682 clknet_1_1__leaf__02672_ VGND VGND VPWR VPWR net714 sky130_fd_sc_hd__inv_2
X_15782_ CPU.registerFile\[13\]\[11\] _03123_ VGND VGND VPWR VPWR _03270_ sky130_fd_sc_hd__or2_1
X_12994_ CPU.registerFile\[5\]\[3\] CPU.registerFile\[4\]\[3\] _04986_ VGND VGND VPWR
+ VPWR _07434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17521_ net710 _01809_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_11945_ _06739_ VGND VGND VPWR VPWR _01598_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17452_ net641 _01740_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[7\] sky130_fd_sc_hd__dfxtp_1
X_11876_ net2466 _05723_ _06697_ VGND VGND VPWR VPWR _06703_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16403_ CPU.registerFile\[16\]\[29\] CPU.registerFile\[18\]\[29\] _05441_ VGND VGND
+ VPWR VPWR _03873_ sky130_fd_sc_hd__mux2_1
X_13615_ CPU.registerFile\[18\]\[21\] CPU.registerFile\[22\]\[21\] _07314_ VGND VGND
+ VPWR VPWR _08037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17383_ net572 _01671_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10827_ _06110_ VGND VGND VPWR VPWR _02090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14595_ clknet_1_0__leaf__07222_ VGND VGND VPWR VPWR _02675_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_119_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16334_ CPU.registerFile\[6\]\[27\] CPU.registerFile\[7\]\[27\] _08395_ VGND VGND
+ VPWR VPWR _03806_ sky130_fd_sc_hd__mux2_1
X_13546_ CPU.registerFile\[8\]\[19\] CPU.registerFile\[12\]\[19\] _07265_ VGND VGND
+ VPWR VPWR _07970_ sky130_fd_sc_hd__mux2_1
X_10758_ _05497_ net1834 _06070_ VGND VGND VPWR VPWR _06074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16265_ CPU.registerFile\[30\]\[25\] CPU.registerFile\[26\]\[25\] _02772_ VGND VGND
+ VPWR VPWR _03739_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13477_ CPU.registerFile\[8\]\[17\] CPU.registerFile\[12\]\[17\] _07638_ VGND VGND
+ VPWR VPWR _07903_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10689_ _06037_ VGND VGND VPWR VPWR _02155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18004_ net1177 _00006_ VGND VGND VPWR VPWR mapped_spi_flash.state\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_132_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14730__830 clknet_1_1__leaf__02689_ VGND VGND VPWR VPWR net862 sky130_fd_sc_hd__inv_2
X_12428_ _05150_ net2419 _07024_ VGND VGND VPWR VPWR _07033_ sky130_fd_sc_hd__mux2_1
X_16196_ CPU.registerFile\[16\]\[23\] CPU.registerFile\[18\]\[23\] _05441_ VGND VGND
+ VPWR VPWR _03672_ sky130_fd_sc_hd__mux2_1
X_12359_ _06996_ VGND VGND VPWR VPWR _01406_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_52_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14648__757 clknet_1_1__leaf__02680_ VGND VGND VPWR VPWR net789 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_147_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_147_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09570_ _04313_ _04701_ VGND VGND VPWR VPWR _05266_ sky130_fd_sc_hd__nor2_1
X_08521_ CPU.aluIn1\[22\] _04239_ VGND VGND VPWR VPWR _04241_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17719_ net908 _02003_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_14935__1015 clknet_1_0__leaf__02709_ VGND VGND VPWR VPWR net1047 sky130_fd_sc_hd__inv_2
XFILLER_0_148_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16658__3 clknet_1_0__leaf__07220_ VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__inv_2
XFILLER_0_156_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14694__799 clknet_1_1__leaf__02684_ VGND VGND VPWR VPWR net831 sky130_fd_sc_hd__inv_2
XFILLER_0_116_611 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14022__301 clknet_1_0__leaf__08362_ VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__inv_2
XFILLER_0_45_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14393__527 clknet_1_0__leaf__02655_ VGND VGND VPWR VPWR net559 sky130_fd_sc_hd__inv_2
X_09004_ CPU.aluIn1\[28\] _04227_ _04699_ VGND VGND VPWR VPWR _04721_ sky130_fd_sc_hd__o21a_1
XFILLER_0_115_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_894 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09906_ _05252_ VGND VGND VPWR VPWR _05539_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_158_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09837_ _05492_ VGND VGND VPWR VPWR _02509_ sky130_fd_sc_hd__clkbuf_1
X_09768_ _05454_ VGND VGND VPWR VPWR _02540_ sky130_fd_sc_hd__clkbuf_1
X_08719_ _04256_ _04331_ VGND VGND VPWR VPWR _04439_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_83_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ _04876_ _05389_ VGND VGND VPWR VPWR _05390_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_83_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ net1311 VGND VGND VPWR VPWR _01694_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11661_ mapped_spi_ram.rcv_data\[28\] _06577_ VGND VGND VPWR VPWR _06582_ sky130_fd_sc_hd__or2_1
X_13400_ CPU.registerFile\[30\]\[14\] CPU.registerFile\[26\]\[14\] _07297_ VGND VGND
+ VPWR VPWR _07829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10612_ net1454 _05981_ VGND VGND VPWR VPWR _05989_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11592_ _06512_ _04635_ VGND VGND VPWR VPWR _06533_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_12_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13331_ CPU.registerFile\[29\]\[12\] _07347_ _07348_ CPU.registerFile\[25\]\[12\]
+ _07349_ VGND VGND VPWR VPWR _07762_ sky130_fd_sc_hd__o221a_1
XFILLER_0_106_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10543_ _05816_ VGND VGND VPWR VPWR _05942_ sky130_fd_sc_hd__clkbuf_4
X_16050_ CPU.aluIn1\[18\] _03081_ _03530_ _03080_ VGND VGND VPWR VPWR _02432_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_114_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13262_ _07474_ _07691_ _07694_ VGND VGND VPWR VPWR _07695_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_114_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10474_ net1377 _05849_ _05884_ _05885_ VGND VGND VPWR VPWR _02217_ sky130_fd_sc_hd__o211a_1
X_12213_ _06859_ VGND VGND VPWR VPWR _06894_ sky130_fd_sc_hd__clkbuf_4
X_13193_ CPU.registerFile\[28\]\[8\] CPU.registerFile\[24\]\[8\] _07399_ VGND VGND
+ VPWR VPWR _07628_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12144_ _05253_ net2226 _06841_ VGND VGND VPWR VPWR _06845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16952_ net247 _01278_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_12075_ _06808_ VGND VGND VPWR VPWR _01536_ sky130_fd_sc_hd__clkbuf_1
X_15903_ CPU.registerFile\[1\]\[14\] _02939_ _03387_ _02943_ VGND VGND VPWR VPWR _03388_
+ sky130_fd_sc_hd__a22o_1
X_11026_ _06216_ VGND VGND VPWR VPWR _01997_ sky130_fd_sc_hd__clkbuf_1
X_16883_ per_uart.uart0.rx_bitcount\[0\] _04164_ _04165_ _05815_ VGND VGND VPWR VPWR
+ _04166_ sky130_fd_sc_hd__a211oi_1
X_15834_ CPU.registerFile\[5\]\[12\] CPU.registerFile\[4\]\[12\] _03146_ VGND VGND
+ VPWR VPWR _03321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15765_ _02851_ VGND VGND VPWR VPWR _03254_ sky130_fd_sc_hd__clkbuf_8
X_12977_ _07417_ VGND VGND VPWR VPWR _07418_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_125_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17504_ net693 _01792_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_11928_ _06730_ VGND VGND VPWR VPWR _01606_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_142_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15696_ CPU.registerFile\[16\]\[8\] _02833_ _02836_ CPU.registerFile\[17\]\[8\] _02764_
+ VGND VGND VPWR VPWR _03187_ sky130_fd_sc_hd__o221a_1
XFILLER_0_86_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17435_ net624 net1461 VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11859_ net2327 _05706_ _06686_ VGND VGND VPWR VPWR _06694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_18 _02887_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17366_ net555 _01654_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[30\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_29 _03064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13529_ CPU.rs2\[18\] _07705_ _07938_ _07953_ _07737_ VGND VGND VPWR VPWR _01313_
+ sky130_fd_sc_hd__o221a_1
X_16317_ _05093_ _03787_ _03788_ _03789_ _03028_ VGND VGND VPWR VPWR _03790_ sky130_fd_sc_hd__o221a_1
X_17297_ net486 _01585_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16248_ CPU.registerFile\[16\]\[24\] _02831_ _02834_ CPU.registerFile\[17\]\[24\]
+ _02854_ VGND VGND VPWR VPWR _03723_ sky130_fd_sc_hd__o221a_1
Xclkbuf_1_1__f__08462_ clknet_0__08462_ VGND VGND VPWR VPWR clknet_1_1__leaf__08462_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16179_ CPU.registerFile\[18\]\[22\] _02833_ _02836_ CPU.registerFile\[19\]\[22\]
+ _03655_ VGND VGND VPWR VPWR _03656_ sky130_fd_sc_hd__o221a_1
XFILLER_0_3_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_149_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09622_ _05286_ _05312_ _05315_ VGND VGND VPWR VPWR _05316_ sky130_fd_sc_hd__and3_1
X_09553_ _05243_ _05249_ _04708_ VGND VGND VPWR VPWR _05250_ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_39_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08504_ CPU.aluIn1\[29\] _04223_ VGND VGND VPWR VPWR _04224_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_65_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09484_ _05182_ _05183_ _04374_ VGND VGND VPWR VPWR _05184_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14401__534 clknet_1_1__leaf__02656_ VGND VGND VPWR VPWR net566 sky130_fd_sc_hd__inv_2
XFILLER_0_58_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15139__1168 clknet_1_0__leaf__02744_ VGND VGND VPWR VPWR net1200 sky130_fd_sc_hd__inv_2
XFILLER_0_61_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10190_ net2321 _05702_ _05692_ VGND VGND VPWR VPWR _05703_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12900_ CPU.registerFile\[13\]\[1\] _07282_ _07341_ VGND VGND VPWR VPWR _07342_ sky130_fd_sc_hd__o21a_1
X_13880_ _07334_ _08283_ _08286_ _08293_ _07766_ VGND VGND VPWR VPWR _08294_ sky130_fd_sc_hd__o311a_1
X_16655__99 clknet_1_1__leaf__03989_ VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__inv_2
X_12831_ _04938_ VGND VGND VPWR VPWR _07274_ sky130_fd_sc_hd__buf_4
XFILLER_0_69_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15550_ _02771_ _03041_ _03042_ _03043_ _02782_ VGND VGND VPWR VPWR _03044_ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11713_ net1330 _06601_ VGND VGND VPWR VPWR _06611_ sky130_fd_sc_hd__or2_1
X_15481_ _08411_ _02967_ _02976_ _08408_ VGND VGND VPWR VPWR _02977_ sky130_fd_sc_hd__o211a_1
X_12693_ _07176_ VGND VGND VPWR VPWR _00038_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17220_ net410 _01508_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_14677__783 clknet_1_1__leaf__02683_ VGND VGND VPWR VPWR net815 sky130_fd_sc_hd__inv_2
X_11644_ _06568_ VGND VGND VPWR VPWR _01727_ sky130_fd_sc_hd__clkbuf_1
X_14376__511 clknet_1_0__leaf__02654_ VGND VGND VPWR VPWR net543 sky130_fd_sc_hd__inv_2
X_17151_ net375 _01439_ VGND VGND VPWR VPWR CPU.aluReg\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11575_ net1361 _06495_ _06521_ _06516_ VGND VGND VPWR VPWR _01749_ sky130_fd_sc_hd__o211a_1
X_16102_ CPU.registerFile\[14\]\[20\] _02889_ VGND VGND VPWR VPWR _03581_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_96_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13314_ CPU.registerFile\[5\]\[12\] CPU.registerFile\[4\]\[12\] _04986_ VGND VGND
+ VPWR VPWR _07745_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17082_ net340 _01404_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_10526_ _05886_ _05929_ VGND VGND VPWR VPWR _05930_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16033_ _02885_ _03511_ _03512_ _03513_ _03054_ VGND VGND VPWR VPWR _03514_ sky130_fd_sc_hd__a221o_1
XFILLER_0_33_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13245_ CPU.registerFile\[3\]\[10\] _07373_ _07376_ VGND VGND VPWR VPWR _07678_ sky130_fd_sc_hd__o21a_1
X_10457_ _04554_ _05869_ _04629_ VGND VGND VPWR VPWR _05871_ sky130_fd_sc_hd__a21o_1
Xclkbuf_1_1__f__02671_ clknet_0__02671_ VGND VGND VPWR VPWR clknet_1_1__leaf__02671_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_149_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14075__349 clknet_1_0__leaf__08367_ VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__inv_2
X_13176_ CPU.registerFile\[1\]\[8\] _07576_ _07610_ _07369_ VGND VGND VPWR VPWR _07611_
+ sky130_fd_sc_hd__a22o_1
X_14934__1014 clknet_1_1__leaf__02709_ VGND VGND VPWR VPWR net1046 sky130_fd_sc_hd__inv_2
X_10388_ mapped_spi_flash.snd_bitcount\[5\] mapped_spi_flash.snd_bitcount\[1\] mapped_spi_flash.snd_bitcount\[0\]
+ mapped_spi_flash.clk_div VGND VGND VPWR VPWR _05818_ sky130_fd_sc_hd__or4bb_1
X_12127_ _05090_ net1899 _06830_ VGND VGND VPWR VPWR _06836_ sky130_fd_sc_hd__mux2_1
X_17984_ net1172 _02268_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_14842__931 clknet_1_1__leaf__02700_ VGND VGND VPWR VPWR net963 sky130_fd_sc_hd__inv_2
X_12058_ _06799_ VGND VGND VPWR VPWR _01544_ sky130_fd_sc_hd__clkbuf_1
X_16935_ clknet_leaf_5_clk _01261_ VGND VGND VPWR VPWR per_uart.uart0.txd_reg\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_127_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11009_ net2388 _05723_ _06201_ VGND VGND VPWR VPWR _06207_ sky130_fd_sc_hd__mux2_1
X_16866_ _03974_ _04152_ _04153_ _04193_ VGND VGND VPWR VPWR _04154_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15817_ CPU.registerFile\[13\]\[12\] _03123_ VGND VGND VPWR VPWR _03304_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16797_ _05288_ _08454_ _04913_ VGND VGND VPWR VPWR _04107_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_36_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15748_ CPU.registerFile\[16\]\[10\] CPU.registerFile\[18\]\[10\] _03032_ VGND VGND
+ VPWR VPWR _03237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_290 _05843_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_15679_ CPU.registerFile\[24\]\[8\] _03130_ _02790_ _03169_ VGND VGND VPWR VPWR _03170_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16567__40 clknet_1_1__leaf__03968_ VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__inv_2
XFILLER_0_157_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17418_ net607 _01706_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_60_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17349_ net538 _01637_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16582__54 clknet_1_0__leaf__03969_ VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__inv_2
XFILLER_0_130_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08984_ _04226_ _04364_ VGND VGND VPWR VPWR _04702_ sky130_fd_sc_hd__xnor2_1
X_09605_ _04672_ _05297_ _05299_ _04768_ VGND VGND VPWR VPWR _05300_ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_0__f__02691_ clknet_0__02691_ VGND VGND VPWR VPWR clknet_1_0__leaf__02691_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09536_ mapped_spi_flash.rcv_data\[16\] _04690_ _04644_ per_uart.rx_avail VGND VGND
+ VPWR VPWR _05233_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09467_ CPU.cycles\[12\] _04503_ _05164_ _04491_ _05167_ VGND VGND VPWR VPWR _05168_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09398_ _04672_ _05101_ VGND VGND VPWR VPWR _05102_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_129_Right_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11360_ _05553_ net2205 _06359_ VGND VGND VPWR VPWR _06393_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15226__136 clknet_1_1__leaf__02753_ VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__inv_2
XFILLER_0_15_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10311_ _04660_ _04661_ VGND VGND VPWR VPWR _05775_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_120_904 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11291_ _06356_ VGND VGND VPWR VPWR _01872_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13030_ CPU.registerFile\[4\]\[4\] _07388_ VGND VGND VPWR VPWR _07469_ sky130_fd_sc_hd__or2_1
X_10242_ _04663_ _04664_ CPU.writeBack _04665_ VGND VGND VPWR VPWR _05738_ sky130_fd_sc_hd__and4b_4
X_14000__281 clknet_1_0__leaf__08360_ VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_91_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10173_ _04981_ VGND VGND VPWR VPWR _05691_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16720_ _08457_ _04040_ _04041_ _04042_ VGND VGND VPWR VPWR _04043_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_109_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13932_ CPU.registerFile\[13\]\[31\] _07361_ _07283_ CPU.registerFile\[9\]\[31\]
+ _07554_ VGND VGND VPWR VPWR _08344_ sky130_fd_sc_hd__o221a_1
XFILLER_0_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13863_ CPU.registerFile\[21\]\[29\] _07347_ _07429_ CPU.registerFile\[17\]\[29\]
+ _07349_ VGND VGND VPWR VPWR _08277_ sky130_fd_sc_hd__o221a_1
XFILLER_0_44_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__08465_ clknet_0__08465_ VGND VGND VPWR VPWR clknet_1_0__leaf__08465_
+ sky130_fd_sc_hd__clkbuf_16
X_12814_ CPU.registerFile\[5\]\[0\] CPU.registerFile\[4\]\[0\] _04986_ VGND VGND VPWR
+ VPWR _07257_ sky130_fd_sc_hd__mux2_1
X_15602_ _02786_ _03092_ _03094_ _02794_ VGND VGND VPWR VPWR _03095_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_122_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13794_ CPU.registerFile\[5\]\[27\] _07577_ _08209_ _07638_ VGND VGND VPWR VPWR _08210_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_122_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18321_ clknet_leaf_15_clk _02601_ VGND VGND VPWR VPWR CPU.PC\[21\] sky130_fd_sc_hd__dfxtp_1
X_15533_ _02763_ VGND VGND VPWR VPWR _03028_ sky130_fd_sc_hd__clkbuf_8
X_12745_ clknet_1_1__leaf__07219_ VGND VGND VPWR VPWR _07220_ sky130_fd_sc_hd__buf_1
XFILLER_0_84_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15464_ CPU.registerFile\[8\]\[3\] CPU.registerFile\[12\]\[3\] _08403_ VGND VGND
+ VPWR VPWR _02960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18252_ net93 _02532_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_12676_ CPU.cycles\[24\] _07164_ VGND VGND VPWR VPWR _07166_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_618 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17203_ net393 _01491_ VGND VGND VPWR VPWR CPU.aluShamt\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11627_ _06556_ VGND VGND VPWR VPWR _01732_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18183_ net214 _02463_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_15395_ CPU.registerFile\[19\]\[1\] CPU.registerFile\[17\]\[1\] _02875_ VGND VGND
+ VPWR VPWR _02893_ sky130_fd_sc_hd__mux2_1
XFILLER_0_154_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17134_ clknet_leaf_26_clk _00038_ VGND VGND VPWR VPWR CPU.cycles\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11558_ _06488_ VGND VGND VPWR VPWR _06508_ sky130_fd_sc_hd__buf_2
XFILLER_0_13_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold608 CPU.registerFile\[26\]\[14\] VGND VGND VPWR VPWR net1849 sky130_fd_sc_hd__dlygate4sd3_1
X_17065_ net323 _01387_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_10509_ _04538_ _04541_ VGND VGND VPWR VPWR _05915_ sky130_fd_sc_hd__and2_1
X_14277_ _08436_ _05289_ _08454_ _08455_ VGND VGND VPWR VPWR _08456_ sky130_fd_sc_hd__a31o_1
Xhold619 CPU.registerFile\[28\]\[12\] VGND VGND VPWR VPWR net1860 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__02723_ clknet_0__02723_ VGND VGND VPWR VPWR clknet_1_1__leaf__02723_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11489_ _05545_ net2247 _06455_ VGND VGND VPWR VPWR _06462_ sky130_fd_sc_hd__mux2_1
X_16016_ CPU.aluIn1\[17\] _02958_ _03478_ _03497_ _02995_ VGND VGND VPWR VPWR _02431_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_110_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13228_ CPU.registerFile\[30\]\[9\] CPU.registerFile\[26\]\[9\] _07492_ VGND VGND
+ VPWR VPWR _07662_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__02754_ _02754_ VGND VGND VPWR VPWR clknet_0__02754_ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f__02654_ clknet_0__02654_ VGND VGND VPWR VPWR clknet_1_1__leaf__02654_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_21_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13159_ CPU.registerFile\[13\]\[7\] _07414_ _07488_ CPU.registerFile\[9\]\[7\] _07489_
+ VGND VGND VPWR VPWR _07595_ sky130_fd_sc_hd__o221a_1
Xclkbuf_0__02685_ _02685_ VGND VGND VPWR VPWR clknet_0__02685_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_20_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14430__560 clknet_1_1__leaf__02659_ VGND VGND VPWR VPWR net592 sky130_fd_sc_hd__inv_2
XFILLER_0_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17967_ net1155 _02251_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_16918_ net1934 _04182_ VGND VGND VPWR VPWR _04188_ sky130_fd_sc_hd__or2_1
X_17898_ net1087 _02182_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15138__1167 clknet_1_1__leaf__02744_ VGND VGND VPWR VPWR net1199 sky130_fd_sc_hd__inv_2
X_16849_ net1552 per_uart.rx_data\[3\] _04139_ VGND VGND VPWR VPWR _04143_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14348__487 clknet_1_1__leaf__08467_ VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13986__269 clknet_1_0__leaf__08358_ VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__inv_2
X_09321_ _05028_ VGND VGND VPWR VPWR _02569_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09252_ _04450_ _04961_ VGND VGND VPWR VPWR _04962_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09183_ _04850_ _04894_ _04848_ VGND VGND VPWR VPWR _04895_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_145_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14058__333 clknet_1_0__leaf__08366_ VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__inv_2
XFILLER_0_101_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14513__635 clknet_1_0__leaf__02667_ VGND VGND VPWR VPWR net667 sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__08428_ clknet_0__08428_ VGND VGND VPWR VPWR clknet_1_1__leaf__08428_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_73_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14251__423 clknet_1_1__leaf__08435_ VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__inv_2
Xclkbuf_1_1__f__08359_ clknet_0__08359_ VGND VGND VPWR VPWR clknet_1_1__leaf__08359_
+ sky130_fd_sc_hd__clkbuf_16
X_08967_ _04367_ _04489_ _04680_ _04685_ VGND VGND VPWR VPWR _04686_ sky130_fd_sc_hd__a211o_1
X_08898_ _04617_ _04614_ VGND VGND VPWR VPWR _04618_ sky130_fd_sc_hd__nor2_4
Xclkbuf_1_0__f__02743_ clknet_0__02743_ VGND VGND VPWR VPWR clknet_1_0__leaf__02743_
+ sky130_fd_sc_hd__clkbuf_16
X_10860_ _06127_ VGND VGND VPWR VPWR _02074_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_104_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_104_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__02674_ clknet_0__02674_ VGND VGND VPWR VPWR clknet_1_0__leaf__02674_
+ sky130_fd_sc_hd__clkbuf_16
X_09519_ _04271_ _04273_ net1288 _04316_ VGND VGND VPWR VPWR _05217_ sky130_fd_sc_hd__a31o_1
X_10791_ _05530_ net1633 _06081_ VGND VGND VPWR VPWR _06091_ sky130_fd_sc_hd__mux2_1
X_14933__1013 clknet_1_1__leaf__02709_ VGND VGND VPWR VPWR net1045 sky130_fd_sc_hd__inv_2
X_12530_ _07087_ VGND VGND VPWR VPWR _01293_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16546__21 clknet_1_1__leaf__03966_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__inv_2
XFILLER_0_53_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12461_ net2182 _05673_ _07049_ VGND VGND VPWR VPWR _07051_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11412_ _06421_ VGND VGND VPWR VPWR _01816_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12392_ _07014_ VGND VGND VPWR VPWR _01391_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16561__35 clknet_1_1__leaf__03967_ VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__inv_2
X_14131_ _08395_ VGND VGND VPWR VPWR _08396_ sky130_fd_sc_hd__clkbuf_4
X_11343_ _06384_ VGND VGND VPWR VPWR _01848_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14789__884 clknet_1_1__leaf__02694_ VGND VGND VPWR VPWR net916 sky130_fd_sc_hd__inv_2
X_11274_ CPU.registerFile\[9\]\[10\] _05715_ _06346_ VGND VGND VPWR VPWR _06348_ sky130_fd_sc_hd__mux2_1
X_14488__612 clknet_1_1__leaf__02665_ VGND VGND VPWR VPWR net644 sky130_fd_sc_hd__inv_2
X_13013_ CPU.registerFile\[29\]\[3\] _07289_ _07290_ CPU.registerFile\[25\]\[3\] _07249_
+ VGND VGND VPWR VPWR _07453_ sky130_fd_sc_hd__o221a_1
X_10225_ _05726_ VGND VGND VPWR VPWR _02323_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17821_ net1010 _02105_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_10156_ net1982 _05679_ _05671_ VGND VGND VPWR VPWR _05680_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17752_ net941 _02036_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10087_ _05640_ VGND VGND VPWR VPWR _02375_ sky130_fd_sc_hd__clkbuf_1
X_16703_ _04027_ _08459_ _05239_ VGND VGND VPWR VPWR _04028_ sky130_fd_sc_hd__a21o_1
X_13915_ CPU.registerFile\[3\]\[31\] _07804_ _07987_ VGND VGND VPWR VPWR _08327_ sky130_fd_sc_hd__o21a_1
X_17683_ net872 _01971_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_14228__403 clknet_1_1__leaf__08432_ VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__inv_2
X_14895_ clknet_1_1__leaf__02697_ VGND VGND VPWR VPWR _02705_ sky130_fd_sc_hd__buf_1
XFILLER_0_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16634_ clknet_1_1__leaf__07219_ VGND VGND VPWR VPWR _03988_ sky130_fd_sc_hd__buf_1
X_13846_ CPU.registerFile\[3\]\[28\] _04986_ _04938_ VGND VGND VPWR VPWR _08261_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13777_ CPU.registerFile\[31\]\[26\] _07402_ _07420_ CPU.registerFile\[27\]\[26\]
+ _07483_ VGND VGND VPWR VPWR _08194_ sky130_fd_sc_hd__o221a_1
X_10989_ _06196_ VGND VGND VPWR VPWR _02014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18304_ clknet_leaf_13_clk _02584_ VGND VGND VPWR VPWR CPU.PC\[4\] sky130_fd_sc_hd__dfxtp_2
X_15516_ _03004_ _03010_ _02879_ VGND VGND VPWR VPWR _03011_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_139_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12728_ _07208_ VGND VGND VPWR VPWR _01257_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_139_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18235_ net76 _02515_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_15447_ CPU.registerFile\[1\]\[2\] _02814_ _02942_ _02943_ VGND VGND VPWR VPWR _02944_
+ sky130_fd_sc_hd__a22o_1
X_12659_ CPU.cycles\[16\] CPU.cycles\[17\] _07154_ VGND VGND VPWR VPWR _07156_ sky130_fd_sc_hd__and3_1
XFILLER_0_127_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18166_ net197 _02446_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_15378_ CPU.registerFile\[2\]\[1\] _02872_ _02873_ CPU.registerFile\[3\]\[1\] _02875_
+ VGND VGND VPWR VPWR _02876_ sky130_fd_sc_hd__a221o_1
X_15209__120 clknet_1_1__leaf__02752_ VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__inv_2
XFILLER_0_20_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_152_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17117_ clknet_leaf_18_clk _00019_ VGND VGND VPWR VPWR CPU.cycles\[13\] sky130_fd_sc_hd__dfxtp_1
Xhold405 CPU.registerFile\[14\]\[12\] VGND VGND VPWR VPWR net1646 sky130_fd_sc_hd__dlygate4sd3_1
X_14329_ clknet_1_0__leaf__08433_ VGND VGND VPWR VPWR _08466_ sky130_fd_sc_hd__buf_1
Xhold416 CPU.registerFile\[11\]\[26\] VGND VGND VPWR VPWR net1657 sky130_fd_sc_hd__dlygate4sd3_1
X_18097_ net160 _02377_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold427 CPU.registerFile\[7\]\[22\] VGND VGND VPWR VPWR net1668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 CPU.registerFile\[4\]\[22\] VGND VGND VPWR VPWR net1679 sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 CPU.registerFile\[14\]\[29\] VGND VGND VPWR VPWR net1690 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__02706_ clknet_0__02706_ VGND VGND VPWR VPWR clknet_1_1__leaf__02706_
+ sky130_fd_sc_hd__clkbuf_16
X_17048_ net306 _01370_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09870_ _05514_ net2089 _05512_ VGND VGND VPWR VPWR _05515_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _04539_ _04540_ VGND VGND VPWR VPWR _04541_ sky130_fd_sc_hd__nor2_1
Xclkbuf_0__02668_ _02668_ VGND VGND VPWR VPWR clknet_0__02668_ sky130_fd_sc_hd__clkbuf_16
Xhold1105 CPU.registerFile\[8\]\[14\] VGND VGND VPWR VPWR net2346 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1116 CPU.registerFile\[12\]\[9\] VGND VGND VPWR VPWR net2357 sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ _04356_ _04469_ _04471_ VGND VGND VPWR VPWR _04472_ sky130_fd_sc_hd__a21oi_1
Xhold1127 CPU.registerFile\[1\]\[17\] VGND VGND VPWR VPWR net2368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1138 CPU.registerFile\[21\]\[23\] VGND VGND VPWR VPWR net2379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1149 CPU.registerFile\[23\]\[3\] VGND VGND VPWR VPWR net2390 sky130_fd_sc_hd__dlygate4sd3_1
X_08683_ _04270_ CPU.aluIn1\[8\] VGND VGND VPWR VPWR _04403_ sky130_fd_sc_hd__and2b_1
X_14701__805 clknet_1_0__leaf__02685_ VGND VGND VPWR VPWR net837 sky130_fd_sc_hd__inv_2
X_15255__162 clknet_1_1__leaf__02756_ VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__inv_2
XFILLER_0_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_138_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09304_ CPU.Jimm\[19\] _04812_ _04989_ CPU.cycles\[19\] VGND VGND VPWR VPWR _05012_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09235_ _04242_ _04452_ _04456_ VGND VGND VPWR VPWR _04946_ sky130_fd_sc_hd__and3_1
XFILLER_0_61_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09166_ _04871_ _04876_ _04877_ VGND VGND VPWR VPWR _04878_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09097_ _04460_ _04682_ VGND VGND VPWR VPWR _04809_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_712 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold950 CPU.registerFile\[19\]\[0\] VGND VGND VPWR VPWR net2191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold961 CPU.registerFile\[20\]\[6\] VGND VGND VPWR VPWR net2202 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold972 CPU.registerFile\[18\]\[7\] VGND VGND VPWR VPWR net2213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold983 per_uart.rx_data\[2\] VGND VGND VPWR VPWR net2224 sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 CPU.registerFile\[1\]\[7\] VGND VGND VPWR VPWR net2235 sky130_fd_sc_hd__dlygate4sd3_1
X_10010_ _05599_ VGND VGND VPWR VPWR _02411_ sky130_fd_sc_hd__clkbuf_1
X_09999_ _05592_ VGND VGND VPWR VPWR _02447_ sky130_fd_sc_hd__clkbuf_1
X_11961_ _06748_ VGND VGND VPWR VPWR _01591_ sky130_fd_sc_hd__clkbuf_1
X_10912_ net1850 _05694_ _06154_ VGND VGND VPWR VPWR _06156_ sky130_fd_sc_hd__mux2_1
X_13700_ CPU.registerFile\[18\]\[24\] CPU.registerFile\[22\]\[24\] _07785_ VGND VGND
+ VPWR VPWR _08119_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_86_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11892_ net2366 _05668_ _06711_ VGND VGND VPWR VPWR _06712_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13969__253 clknet_1_0__leaf__08357_ VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__inv_2
XFILLER_0_79_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13631_ CPU.registerFile\[3\]\[22\] _07804_ _07987_ VGND VGND VPWR VPWR _08052_ sky130_fd_sc_hd__o21a_1
X_10843_ net1936 _05694_ _06117_ VGND VGND VPWR VPWR _06119_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_0__f__02657_ clknet_0__02657_ VGND VGND VPWR VPWR clknet_1_0__leaf__02657_
+ sky130_fd_sc_hd__clkbuf_16
X_13562_ CPU.registerFile\[6\]\[20\] CPU.registerFile\[7\]\[20\] _07641_ VGND VGND
+ VPWR VPWR _07985_ sky130_fd_sc_hd__mux2_1
X_16350_ _02758_ _03819_ _03821_ _08396_ VGND VGND VPWR VPWR _03822_ sky130_fd_sc_hd__a211o_1
X_10774_ _06082_ VGND VGND VPWR VPWR _02115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12513_ net2061 _05725_ _07071_ VGND VGND VPWR VPWR _07078_ sky130_fd_sc_hd__mux2_1
X_15301_ _02760_ VGND VGND VPWR VPWR _02800_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16281_ _03749_ _03754_ _05361_ VGND VGND VPWR VPWR _03755_ sky130_fd_sc_hd__o21a_1
XFILLER_0_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13493_ CPU.registerFile\[1\]\[17\] _07255_ _07918_ _07638_ VGND VGND VPWR VPWR _07919_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14223__399 clknet_1_0__leaf__08431_ VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__inv_2
X_18020_ net1193 _02300_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_12444_ _07041_ VGND VGND VPWR VPWR _01366_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15163_ clknet_1_0__leaf__02720_ VGND VGND VPWR VPWR _02747_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_117_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_829 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12375_ _05306_ net1935 _06999_ VGND VGND VPWR VPWR _07005_ sky130_fd_sc_hd__mux2_1
X_15137__1166 clknet_1_1__leaf__02744_ VGND VGND VPWR VPWR net1198 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_134_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14114_ _08385_ VGND VGND VPWR VPWR _01466_ sky130_fd_sc_hd__clkbuf_1
X_11326_ _06375_ VGND VGND VPWR VPWR _01856_ sky130_fd_sc_hd__clkbuf_1
X_15094_ net1466 _07185_ VGND VGND VPWR VPWR _02734_ sky130_fd_sc_hd__nand2_1
X_11257_ CPU.registerFile\[9\]\[18\] _05698_ _06335_ VGND VGND VPWR VPWR _06339_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_130_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10208_ _05208_ VGND VGND VPWR VPWR _05715_ sky130_fd_sc_hd__clkbuf_4
X_11188_ _06302_ VGND VGND VPWR VPWR _01921_ sky130_fd_sc_hd__clkbuf_1
X_17804_ net993 _02088_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_10139_ _05667_ VGND VGND VPWR VPWR _02350_ sky130_fd_sc_hd__clkbuf_1
X_15996_ _03252_ _03469_ _03477_ _02935_ VGND VGND VPWR VPWR _03478_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_50_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17735_ net924 _02019_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_17666_ net855 _01954_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_14542__661 clknet_1_0__leaf__02670_ VGND VGND VPWR VPWR net693 sky130_fd_sc_hd__inv_2
X_16617_ net1591 net1565 _03979_ VGND VGND VPWR VPWR _03984_ sky130_fd_sc_hd__mux2_1
X_13829_ CPU.registerFile\[29\]\[28\] _07772_ _07773_ CPU.registerFile\[25\]\[28\]
+ _08243_ VGND VGND VPWR VPWR _08244_ sky130_fd_sc_hd__o221a_1
X_17597_ net786 _01885_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16479_ CPU.registerFile\[15\]\[31\] CPU.registerFile\[11\]\[31\] _02849_ VGND VGND
+ VPWR VPWR _03947_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09020_ _04359_ _04735_ VGND VGND VPWR VPWR _04736_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18218_ net59 _02498_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14198__376 clknet_1_1__leaf__08429_ VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__inv_2
XFILLER_0_142_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18149_ clknet_leaf_26_clk _02429_ VGND VGND VPWR VPWR CPU.aluIn1\[15\] sky130_fd_sc_hd__dfxtp_4
Xhold202 mapped_spi_flash.rcv_data\[22\] VGND VGND VPWR VPWR net1443 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold213 mapped_spi_flash.rcv_data\[16\] VGND VGND VPWR VPWR net1454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 per_uart.uart0.enable16_counter\[13\] VGND VGND VPWR VPWR net1465 sky130_fd_sc_hd__dlygate4sd3_1
X_16540__16 clknet_1_1__leaf__03965_ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__inv_2
Xhold235 mapped_spi_flash.rcv_data\[27\] VGND VGND VPWR VPWR net1476 sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 CPU.cycles\[14\] VGND VGND VPWR VPWR net1487 sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 CPU.state\[0\] VGND VGND VPWR VPWR net1498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 _04140_ VGND VGND VPWR VPWR net1509 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09922_ _05549_ net2059 _05533_ VGND VGND VPWR VPWR _05550_ sky130_fd_sc_hd__mux2_1
Xhold279 _04173_ VGND VGND VPWR VPWR net1520 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14932__1012 clknet_1_0__leaf__02709_ VGND VGND VPWR VPWR net1044 sky130_fd_sc_hd__inv_2
X_09853_ _04779_ VGND VGND VPWR VPWR _05503_ sky130_fd_sc_hd__buf_2
X_08804_ CPU.aluIn1\[0\] _04523_ VGND VGND VPWR VPWR _04524_ sky130_fd_sc_hd__nand2_4
X_09784_ _05462_ VGND VGND VPWR VPWR _02532_ sky130_fd_sc_hd__clkbuf_1
X_14625__736 clknet_1_1__leaf__02678_ VGND VGND VPWR VPWR net768 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_29_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08735_ CPU.aluIn1\[20\] _04454_ _04450_ VGND VGND VPWR VPWR _04455_ sky130_fd_sc_hd__and3_1
XANTENNA_108 _05406_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_08666_ CPU.aluIn1\[18\] VGND VGND VPWR VPWR _04386_ sky130_fd_sc_hd__inv_2
XANTENNA_119 _05516_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08597_ CPU.aluIn1\[9\] _04268_ VGND VGND VPWR VPWR _04317_ sky130_fd_sc_hd__and2_1
XFILLER_0_119_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09218_ CPU.PC\[23\] _04929_ VGND VGND VPWR VPWR _04930_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10490_ _04546_ _05898_ _04629_ VGND VGND VPWR VPWR _05899_ sky130_fd_sc_hd__a21oi_1
X_14671__778 clknet_1_0__leaf__02682_ VGND VGND VPWR VPWR net810 sky130_fd_sc_hd__inv_2
X_09149_ CPU.Bimm\[7\] _04819_ CPU.PC\[7\] VGND VGND VPWR VPWR _04861_ sky130_fd_sc_hd__a21o_1
XFILLER_0_133_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12160_ _05448_ net2021 _06818_ VGND VGND VPWR VPWR _06853_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11111_ _06261_ VGND VGND VPWR VPWR _01957_ sky130_fd_sc_hd__clkbuf_1
X_12091_ _06816_ VGND VGND VPWR VPWR _01528_ sky130_fd_sc_hd__clkbuf_1
Xhold780 CPU.registerFile\[27\]\[0\] VGND VGND VPWR VPWR net2021 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold791 CPU.registerFile\[1\]\[25\] VGND VGND VPWR VPWR net2032 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11042_ _06224_ VGND VGND VPWR VPWR _01989_ sky130_fd_sc_hd__clkbuf_1
X_15850_ _02759_ _03333_ _03335_ _02767_ VGND VGND VPWR VPWR _03336_ sky130_fd_sc_hd__a211o_1
X_15781_ CPU.registerFile\[15\]\[11\] CPU.registerFile\[11\]\[11\] _02773_ VGND VGND
+ VPWR VPWR _03269_ sky130_fd_sc_hd__mux2_1
X_12993_ _07428_ _07432_ _07320_ VGND VGND VPWR VPWR _07433_ sky130_fd_sc_hd__mux2_2
X_17520_ net709 _01808_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_11944_ CPU.registerFile\[11\]\[6\] _05723_ _06733_ VGND VGND VPWR VPWR _06739_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17451_ net640 _01739_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[6\] sky130_fd_sc_hd__dfxtp_1
X_11875_ _06702_ VGND VGND VPWR VPWR _01631_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__02709_ clknet_0__02709_ VGND VGND VPWR VPWR clknet_1_0__leaf__02709_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_129_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16402_ _03022_ _03869_ _03870_ _03871_ _03028_ VGND VGND VPWR VPWR _03872_ sky130_fd_sc_hd__o221a_1
X_10826_ net1881 _05677_ _06106_ VGND VGND VPWR VPWR _06110_ sky130_fd_sc_hd__mux2_1
X_13614_ _07519_ _08034_ _08035_ VGND VGND VPWR VPWR _08036_ sky130_fd_sc_hd__o21ai_1
X_17382_ net571 _01670_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_119_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16333_ CPU.registerFile\[1\]\[27\] _02873_ _03804_ _08404_ VGND VGND VPWR VPWR _03805_
+ sky130_fd_sc_hd__a22o_1
X_13545_ _07961_ _07968_ _07395_ VGND VGND VPWR VPWR _07969_ sky130_fd_sc_hd__o21a_1
X_10757_ _06073_ VGND VGND VPWR VPWR _02123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13476_ _07653_ _07900_ _07901_ VGND VGND VPWR VPWR _07902_ sky130_fd_sc_hd__o21a_1
X_16264_ _02812_ _03735_ _03737_ _02965_ VGND VGND VPWR VPWR _03738_ sky130_fd_sc_hd__a211o_1
XFILLER_0_54_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10688_ _05495_ net1650 _06034_ VGND VGND VPWR VPWR _06037_ sky130_fd_sc_hd__mux2_1
X_18003_ net1176 _00005_ VGND VGND VPWR VPWR mapped_spi_flash.state\[1\] sky130_fd_sc_hd__dfxtp_1
X_12427_ _07032_ VGND VGND VPWR VPWR _01374_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_132_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16195_ _02885_ _03667_ _03668_ _03670_ VGND VGND VPWR VPWR _03671_ sky130_fd_sc_hd__o22a_1
X_12358_ _05130_ net2043 _06988_ VGND VGND VPWR VPWR _06996_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11309_ _06366_ VGND VGND VPWR VPWR _01864_ sky130_fd_sc_hd__clkbuf_1
X_12289_ CPU.aluReg\[8\] CPU.aluReg\[6\] _06939_ VGND VGND VPWR VPWR _06952_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_147_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15979_ _02936_ _03454_ _03461_ _02934_ VGND VGND VPWR VPWR _03462_ sky130_fd_sc_hd__o211a_1
X_08520_ CPU.aluIn1\[22\] _04239_ VGND VGND VPWR VPWR _04240_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15029__1100 clknet_1_1__leaf__02718_ VGND VGND VPWR VPWR net1132 sky130_fd_sc_hd__inv_2
X_17718_ net907 _02002_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17649_ net838 _01937_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_11_Left_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14206__383 clknet_1_0__leaf__08430_ VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__inv_2
X_14813__906 clknet_1_0__leaf__02696_ VGND VGND VPWR VPWR net938 sky130_fd_sc_hd__inv_2
XFILLER_0_116_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09003_ CPU.Bimm\[8\] _04498_ _04503_ CPU.cycles\[28\] _04719_ VGND VGND VPWR VPWR
+ _04720_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12753__206 clknet_1_1__leaf__07221_ VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__inv_2
XFILLER_0_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09905_ _05538_ VGND VGND VPWR VPWR _02487_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09836_ _05487_ net2272 _05491_ VGND VGND VPWR VPWR _05492_ sky130_fd_sc_hd__mux2_1
X_09767_ net1743 _04696_ _05452_ VGND VGND VPWR VPWR _05454_ sky130_fd_sc_hd__mux2_1
X_08718_ _04396_ _04436_ _04437_ VGND VGND VPWR VPWR _04438_ sky130_fd_sc_hd__o21a_1
XFILLER_0_69_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09698_ CPU.PC\[1\] _04872_ _04875_ VGND VGND VPWR VPWR _05389_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_83_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15136__1165 clknet_1_1__leaf__02744_ VGND VGND VPWR VPWR net1197 sky130_fd_sc_hd__inv_2
XFILLER_0_68_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ CPU.aluIn1\[31\] VGND VGND VPWR VPWR _04369_ sky130_fd_sc_hd__inv_2
XFILLER_0_139_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11660_ net1463 _06575_ _06580_ _06581_ VGND VGND VPWR VPWR _01724_ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10611_ net1454 _05983_ _05988_ _05980_ VGND VGND VPWR VPWR _02183_ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11591_ net1375 _06524_ _06532_ _06516_ VGND VGND VPWR VPWR _01744_ sky130_fd_sc_hd__o211a_1
XFILLER_0_119_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13330_ CPU.registerFile\[31\]\[12\] _07556_ _07557_ CPU.registerFile\[27\]\[12\]
+ _07345_ VGND VGND VPWR VPWR _07761_ sky130_fd_sc_hd__o221a_1
XFILLER_0_107_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10542_ _05813_ _05821_ net1528 VGND VGND VPWR VPWR _05941_ sky130_fd_sc_hd__o21a_1
XFILLER_0_51_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13261_ CPU.registerFile\[27\]\[10\] _07363_ _07693_ VGND VGND VPWR VPWR _07694_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_98_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10473_ _05843_ VGND VGND VPWR VPWR _05885_ sky130_fd_sc_hd__buf_2
XFILLER_0_134_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12212_ CPU.aluReg\[26\] CPU.aluReg\[24\] _06871_ VGND VGND VPWR VPWR _06893_ sky130_fd_sc_hd__mux2_1
X_13192_ _07411_ _07623_ _07626_ VGND VGND VPWR VPWR _07627_ sky130_fd_sc_hd__or3_1
XFILLER_0_103_873 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12143_ _06844_ VGND VGND VPWR VPWR _01504_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16951_ net246 _01277_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_12074_ _05230_ net1957 _06805_ VGND VGND VPWR VPWR _06808_ sky130_fd_sc_hd__mux2_1
X_14909__992 clknet_1_1__leaf__02706_ VGND VGND VPWR VPWR net1024 sky130_fd_sc_hd__inv_2
X_15195__108 clknet_1_0__leaf__02750_ VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__inv_2
X_15902_ CPU.registerFile\[5\]\[14\] CPU.registerFile\[4\]\[14\] _03146_ VGND VGND
+ VPWR VPWR _03387_ sky130_fd_sc_hd__mux2_1
X_11025_ net1739 _05668_ _06215_ VGND VGND VPWR VPWR _06216_ sky130_fd_sc_hd__mux2_1
X_16882_ _03972_ _04151_ _08355_ VGND VGND VPWR VPWR _04165_ sky130_fd_sc_hd__and3_1
X_14608__720 clknet_1_0__leaf__02677_ VGND VGND VPWR VPWR net752 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_129_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15833_ CPU.registerFile\[2\]\[12\] _03143_ _02980_ CPU.registerFile\[3\]\[12\] _03144_
+ VGND VGND VPWR VPWR _03320_ sky130_fd_sc_hd__a221o_1
XFILLER_0_154_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15764_ _03246_ _03251_ _03252_ VGND VGND VPWR VPWR _03253_ sky130_fd_sc_hd__a21o_1
X_12976_ _05338_ VGND VGND VPWR VPWR _07417_ sky130_fd_sc_hd__clkbuf_8
X_17503_ net692 _01791_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_142_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11927_ CPU.registerFile\[11\]\[14\] _05706_ _06722_ VGND VGND VPWR VPWR _06730_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_142_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15695_ CPU.registerFile\[20\]\[8\] CPU.registerFile\[21\]\[8\] _08395_ VGND VGND
+ VPWR VPWR _03186_ sky130_fd_sc_hd__mux2_1
X_17434_ net623 net1413 VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[27\] sky130_fd_sc_hd__dfxtp_1
X_11858_ _06693_ VGND VGND VPWR VPWR _01639_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14931__1011 clknet_1_1__leaf__02709_ VGND VGND VPWR VPWR net1043 sky130_fd_sc_hd__inv_2
XFILLER_0_28_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17365_ net554 _01653_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[29\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_19 _02895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_10809_ _06100_ VGND VGND VPWR VPWR _02098_ sky130_fd_sc_hd__clkbuf_1
X_11789_ _05109_ net2534 _06650_ VGND VGND VPWR VPWR _06657_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_126_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16316_ CPU.registerFile\[20\]\[26\] _03025_ _02829_ VGND VGND VPWR VPWR _03789_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13528_ _07306_ _07945_ _07952_ _07703_ VGND VGND VPWR VPWR _07953_ sky130_fd_sc_hd__a31o_1
X_17296_ net485 _01584_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14654__762 clknet_1_1__leaf__02681_ VGND VGND VPWR VPWR net794 sky130_fd_sc_hd__inv_2
XFILLER_0_152_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16247_ CPU.registerFile\[20\]\[24\] CPU.registerFile\[21\]\[24\] _08394_ VGND VGND
+ VPWR VPWR _03722_ sky130_fd_sc_hd__mux2_1
X_13459_ CPU.registerFile\[8\]\[16\] CPU.registerFile\[12\]\[16\] _05283_ VGND VGND
+ VPWR VPWR _07886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_152_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16178_ _03065_ _03654_ VGND VGND VPWR VPWR _03655_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16925__5 clknet_1_1__leaf__07220_ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_149_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14052__328 clknet_1_1__leaf__08365_ VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__inv_2
XFILLER_0_128_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09621_ _05275_ _05133_ _05314_ _04484_ VGND VGND VPWR VPWR _05315_ sky130_fd_sc_hd__o22a_1
X_09552_ _04426_ _04806_ _05248_ _04679_ VGND VGND VPWR VPWR _05249_ sky130_fd_sc_hd__a2bb2o_1
X_08503_ CPU.rs2\[29\] _04201_ _04206_ VGND VGND VPWR VPWR _04223_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_65_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09483_ _04323_ _05159_ VGND VGND VPWR VPWR _05183_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14737__837 clknet_1_0__leaf__02689_ VGND VGND VPWR VPWR net869 sky130_fd_sc_hd__inv_2
XFILLER_0_58_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_784 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15052__1119 clknet_1_0__leaf__02721_ VGND VGND VPWR VPWR net1151 sky130_fd_sc_hd__inv_2
XFILLER_0_14_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14783__879 clknet_1_0__leaf__02693_ VGND VGND VPWR VPWR net911 sky130_fd_sc_hd__inv_2
X_09819_ net2165 _05333_ _05474_ VGND VGND VPWR VPWR _05481_ sky130_fd_sc_hd__mux2_1
X_12830_ _07272_ VGND VGND VPWR VPWR _07273_ sky130_fd_sc_hd__buf_4
XFILLER_0_68_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_158_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14029__308 clknet_1_0__leaf__08362_ VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__inv_2
XFILLER_0_57_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11712_ net1330 _06603_ _06610_ _06607_ VGND VGND VPWR VPWR _01701_ sky130_fd_sc_hd__o211a_1
X_12692_ _07174_ _07175_ VGND VGND VPWR VPWR _07176_ sky130_fd_sc_hd__and2_1
X_15480_ _02971_ _02975_ _02879_ VGND VGND VPWR VPWR _02976_ sky130_fd_sc_hd__a21o_1
X_11643_ _06492_ _06562_ mapped_spi_ram.snd_bitcount\[0\] VGND VGND VPWR VPWR _06568_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17150_ net374 _01438_ VGND VGND VPWR VPWR CPU.aluReg\[14\] sky130_fd_sc_hd__dfxtp_1
X_14362_ clknet_1_0__leaf__08433_ VGND VGND VPWR VPWR _02652_ sky130_fd_sc_hd__buf_1
X_11574_ net1371 _06517_ _06509_ _06520_ VGND VGND VPWR VPWR _06521_ sky130_fd_sc_hd__a211o_1
XFILLER_0_25_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16101_ CPU.registerFile\[8\]\[20\] CPU.registerFile\[12\]\[20\] _03254_ VGND VGND
+ VPWR VPWR _03580_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10525_ CPU.PC\[5\] _04598_ _05927_ _05928_ VGND VGND VPWR VPWR _05929_ sky130_fd_sc_hd__o2bb2a_1
X_13313_ _07740_ _07743_ _07320_ VGND VGND VPWR VPWR _07744_ sky130_fd_sc_hd__mux2_4
XFILLER_0_52_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17081_ net339 _01403_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_13244_ CPU.registerFile\[2\]\[10\] _07322_ VGND VGND VPWR VPWR _07677_ sky130_fd_sc_hd__or2_1
X_16032_ CPU.registerFile\[25\]\[18\] _03280_ _02940_ VGND VGND VPWR VPWR _03513_
+ sky130_fd_sc_hd__o21a_1
X_10456_ _04554_ _05869_ VGND VGND VPWR VPWR _05870_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__02670_ clknet_0__02670_ VGND VGND VPWR VPWR clknet_1_1__leaf__02670_
+ sky130_fd_sc_hd__clkbuf_16
X_13175_ CPU.registerFile\[5\]\[8\] CPU.registerFile\[4\]\[8\] _07577_ VGND VGND VPWR
+ VPWR _07610_ sky130_fd_sc_hd__mux2_1
X_15203__115 clknet_1_0__leaf__02751_ VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__inv_2
X_10387_ mapped_spi_flash.state\[1\] VGND VGND VPWR VPWR _05817_ sky130_fd_sc_hd__clkbuf_2
X_12126_ _06835_ VGND VGND VPWR VPWR _01512_ sky130_fd_sc_hd__clkbuf_1
X_17983_ net1171 _02267_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[28\] sky130_fd_sc_hd__dfxtp_1
X_12057_ net1244 net2201 _06794_ VGND VGND VPWR VPWR _06799_ sky130_fd_sc_hd__mux2_1
X_16934_ clknet_leaf_7_clk _01260_ VGND VGND VPWR VPWR per_uart.uart0.txd_reg\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_144_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11008_ _06206_ VGND VGND VPWR VPWR _02005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_144_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16865_ _03972_ per_uart.uart0.uart_rxd2 _07195_ VGND VGND VPWR VPWR _04153_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_88_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15816_ CPU.registerFile\[15\]\[12\] CPU.registerFile\[11\]\[12\] _02773_ VGND VGND
+ VPWR VPWR _03303_ sky130_fd_sc_hd__mux2_1
X_16796_ net1762 _04032_ VGND VGND VPWR VPWR _04106_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_36_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15747_ _03022_ _03233_ _03234_ _03235_ _02895_ VGND VGND VPWR VPWR _03236_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_47_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12959_ CPU.registerFile\[30\]\[2\] CPU.registerFile\[26\]\[2\] _07399_ VGND VGND
+ VPWR VPWR _07400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15678_ CPU.registerFile\[28\]\[8\] _02791_ VGND VGND VPWR VPWR _03169_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_280 _05551_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_291 _07084_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17417_ net606 _01705_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[10\] sky130_fd_sc_hd__dfxtp_1
X_14629_ clknet_1_0__leaf__02675_ VGND VGND VPWR VPWR _02679_ sky130_fd_sc_hd__buf_1
XFILLER_0_23_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17348_ net537 _01636_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17279_ net468 _01567_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15135__1164 clknet_1_1__leaf__02744_ VGND VGND VPWR VPWR net1196 sky130_fd_sc_hd__inv_2
XFILLER_0_2_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_58_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08983_ CPU.Jimm\[14\] _04487_ VGND VGND VPWR VPWR _04701_ sky130_fd_sc_hd__nand2_4
XFILLER_0_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09604_ _04800_ _05298_ VGND VGND VPWR VPWR _05299_ sky130_fd_sc_hd__nand2_1
XFILLER_0_97_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__02690_ clknet_0__02690_ VGND VGND VPWR VPWR clknet_1_0__leaf__02690_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09535_ mapped_spi_ram.rcv_data\[0\] _04688_ _04709_ mapped_spi_flash.rcv_data\[0\]
+ VGND VGND VPWR VPWR _05232_ sky130_fd_sc_hd__a22o_4
X_09466_ _04818_ _05166_ VGND VGND VPWR VPWR _05167_ sky130_fd_sc_hd__nor2_1
X_14325__466 clknet_1_0__leaf__08465_ VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__inv_2
XFILLER_0_149_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09397_ _04330_ _04439_ VGND VGND VPWR VPWR _05101_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_136_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_468 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13963__248 clknet_1_1__leaf__08356_ VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__inv_2
XFILLER_0_74_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_913 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10310_ _05774_ VGND VGND VPWR VPWR _02286_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11290_ CPU.registerFile\[9\]\[2\] _05731_ _06346_ VGND VGND VPWR VPWR _06356_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10241_ _04660_ _04661_ VGND VGND VPWR VPWR _05737_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_91_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10172_ _05690_ VGND VGND VPWR VPWR _02340_ sky130_fd_sc_hd__clkbuf_1
X_14035__312 clknet_1_0__leaf__08364_ VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__inv_2
XFILLER_0_100_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14930__1010 clknet_1_1__leaf__02709_ VGND VGND VPWR VPWR net1042 sky130_fd_sc_hd__inv_2
X_12766__216 clknet_1_0__leaf__07224_ VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_109_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13931_ CPU.registerFile\[8\]\[31\] CPU.registerFile\[12\]\[31\] _07785_ VGND VGND
+ VPWR VPWR _08343_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_109_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13862_ CPU.registerFile\[16\]\[29\] CPU.registerFile\[20\]\[29\] _07648_ VGND VGND
+ VPWR VPWR _08276_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__08464_ clknet_0__08464_ VGND VGND VPWR VPWR clknet_1_0__leaf__08464_
+ sky130_fd_sc_hd__clkbuf_16
X_15601_ CPU.registerFile\[24\]\[6\] _02789_ _02790_ _03093_ VGND VGND VPWR VPWR _03094_
+ sky130_fd_sc_hd__o211a_1
X_12813_ _07255_ VGND VGND VPWR VPWR _07256_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_2_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_122_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13793_ CPU.registerFile\[4\]\[27\] _07374_ VGND VGND VPWR VPWR _08209_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_122_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18320_ clknet_leaf_15_clk _02600_ VGND VGND VPWR VPWR CPU.PC\[20\] sky130_fd_sc_hd__dfxtp_1
X_15532_ CPU.registerFile\[20\]\[4\] _03025_ _03026_ VGND VGND VPWR VPWR _03027_ sky130_fd_sc_hd__a21o_1
X_12744_ clknet_leaf_0_clk VGND VGND VPWR VPWR _07219_ sky130_fd_sc_hd__buf_1
X_18251_ net92 _02531_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_15463_ CPU.registerFile\[14\]\[3\] CPU.registerFile\[10\]\[3\] _02906_ VGND VGND
+ VPWR VPWR _02959_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14081__354 clknet_1_0__leaf__08368_ VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__inv_2
X_12675_ _07164_ net1438 VGND VGND VPWR VPWR _00030_ sky130_fd_sc_hd__nor2_1
X_17202_ net392 _01490_ VGND VGND VPWR VPWR CPU.aluShamt\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_42_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18182_ net213 _02462_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_42_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11626_ net2439 _06554_ _06555_ VGND VGND VPWR VPWR _06556_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_693 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15394_ _02848_ _02884_ _02891_ _02843_ VGND VGND VPWR VPWR _02892_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_100_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17133_ clknet_leaf_22_clk _00036_ VGND VGND VPWR VPWR CPU.cycles\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_663 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11557_ net1389 _06495_ _06507_ _06006_ VGND VGND VPWR VPWR _01753_ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold609 CPU.registerFile\[5\]\[20\] VGND VGND VPWR VPWR net1850 sky130_fd_sc_hd__dlygate4sd3_1
X_17064_ net322 _01386_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_10508_ CPU.aluIn1\[7\] CPU.Bimm\[7\] VGND VGND VPWR VPWR _05914_ sky130_fd_sc_hd__nand2_1
Xclkbuf_1_1__f__02722_ clknet_0__02722_ VGND VGND VPWR VPWR clknet_1_1__leaf__02722_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14276_ CPU.state\[1\] VGND VGND VPWR VPWR _08455_ sky130_fd_sc_hd__inv_2
X_11488_ _06461_ VGND VGND VPWR VPWR _01780_ sky130_fd_sc_hd__clkbuf_1
X_16015_ _08408_ _03487_ _03496_ _02993_ VGND VGND VPWR VPWR _03497_ sky130_fd_sc_hd__a31o_1
X_13227_ _07412_ _07659_ _07660_ VGND VGND VPWR VPWR _07661_ sky130_fd_sc_hd__o21a_1
X_10439_ _05856_ _05857_ VGND VGND VPWR VPWR _05858_ sky130_fd_sc_hd__or2_1
Xclkbuf_0__02753_ _02753_ VGND VGND VPWR VPWR clknet_0__02753_ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f__02653_ clknet_0__02653_ VGND VGND VPWR VPWR clknet_1_1__leaf__02653_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_21_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13158_ CPU.registerFile\[8\]\[7\] CPU.registerFile\[12\]\[7\] _07265_ VGND VGND
+ VPWR VPWR _07594_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__02684_ _02684_ VGND VGND VPWR VPWR clknet_0__02684_ sky130_fd_sc_hd__clkbuf_16
X_14766__863 clknet_1_0__leaf__02692_ VGND VGND VPWR VPWR net895 sky130_fd_sc_hd__inv_2
X_12109_ _06826_ VGND VGND VPWR VPWR _01520_ sky130_fd_sc_hd__clkbuf_1
X_13089_ CPU.registerFile\[29\]\[5\] _07347_ _07348_ CPU.registerFile\[25\]\[5\] _07349_
+ VGND VGND VPWR VPWR _07527_ sky130_fd_sc_hd__o221a_1
X_17966_ net1154 _02250_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_16526__193 clknet_1_0__leaf__03964_ VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__inv_2
XFILLER_0_18_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16917_ CPU.mem_wdata\[4\] _04180_ _04187_ _04176_ VGND VGND VPWR VPWR _02642_ sky130_fd_sc_hd__o211a_1
X_17897_ net1086 _02181_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[15\] sky130_fd_sc_hd__dfxtp_1
X_16848_ _04142_ VGND VGND VPWR VPWR _02618_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16779_ _04027_ _04039_ _05003_ VGND VGND VPWR VPWR _04092_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15051__1118 clknet_1_0__leaf__02721_ VGND VGND VPWR VPWR net1150 sky130_fd_sc_hd__inv_2
XFILLER_0_76_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09320_ net1559 _05027_ _04983_ VGND VGND VPWR VPWR _05028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09251_ CPU.aluIn1\[20\] _04454_ _04960_ VGND VGND VPWR VPWR _04961_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_157_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_157_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09182_ _04852_ _04892_ _04893_ VGND VGND VPWR VPWR _04894_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_888 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03969_ clknet_0__03969_ VGND VGND VPWR VPWR clknet_1_1__leaf__03969_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14849__938 clknet_1_0__leaf__02700_ VGND VGND VPWR VPWR net970 sky130_fd_sc_hd__inv_2
XFILLER_0_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__08358_ clknet_0__08358_ VGND VGND VPWR VPWR clknet_1_1__leaf__08358_
+ sky130_fd_sc_hd__clkbuf_16
X_08966_ _04366_ _04211_ _04681_ CPU.aluReg\[30\] _04684_ VGND VGND VPWR VPWR _04685_
+ sky130_fd_sc_hd__a221o_1
X_08897_ _04611_ _04615_ _04616_ _04608_ VGND VGND VPWR VPWR _04617_ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_3_Left_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_0__f__02673_ clknet_0__02673_ VGND VGND VPWR VPWR clknet_1_0__leaf__02673_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_104_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09518_ _04429_ _05215_ VGND VGND VPWR VPWR _05216_ sky130_fd_sc_hd__nor2_1
X_10790_ _06090_ VGND VGND VPWR VPWR _02107_ sky130_fd_sc_hd__clkbuf_1
X_15232__141 clknet_1_1__leaf__02754_ VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__inv_2
XFILLER_0_137_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09449_ CPU.registerFile\[16\]\[13\] _05150_ _04983_ VGND VGND VPWR VPWR _05151_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_811 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12460_ _07050_ VGND VGND VPWR VPWR _01359_ sky130_fd_sc_hd__clkbuf_1
X_11411_ _05535_ CPU.registerFile\[24\]\[10\] _06419_ VGND VGND VPWR VPWR _06421_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12391_ _04659_ net1962 _07013_ VGND VGND VPWR VPWR _07014_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11342_ _05535_ CPU.registerFile\[23\]\[10\] _06382_ VGND VGND VPWR VPWR _06384_
+ sky130_fd_sc_hd__mux2_1
X_14130_ _08394_ VGND VGND VPWR VPWR _08395_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_105_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11273_ _06347_ VGND VGND VPWR VPWR _01881_ sky130_fd_sc_hd__clkbuf_1
X_10224_ net1724 _05725_ _05713_ VGND VGND VPWR VPWR _05726_ sky130_fd_sc_hd__mux2_1
X_13012_ _07296_ _07451_ VGND VGND VPWR VPWR _07452_ sky130_fd_sc_hd__or2_1
X_17820_ net1009 _02104_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10155_ _04747_ VGND VGND VPWR VPWR _05679_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_7_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17751_ net940 _02035_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_10086_ net1671 _04780_ _05633_ VGND VGND VPWR VPWR _05640_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16702_ _05288_ VGND VGND VPWR VPWR _04027_ sky130_fd_sc_hd__buf_2
X_13914_ CPU.registerFile\[2\]\[31\] _07621_ VGND VGND VPWR VPWR _08326_ sky130_fd_sc_hd__or2_1
Xclkbuf_1_0__f__03989_ clknet_0__03989_ VGND VGND VPWR VPWR clknet_1_0__leaf__03989_
+ sky130_fd_sc_hd__clkbuf_16
X_17682_ net871 _01970_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_13845_ CPU.registerFile\[2\]\[28\] _07388_ VGND VGND VPWR VPWR _08260_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14308__450 clknet_1_0__leaf__08464_ VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__inv_2
X_15134__1163 clknet_1_1__leaf__02744_ VGND VGND VPWR VPWR net1195 sky130_fd_sc_hd__inv_2
X_13776_ CPU.registerFile\[30\]\[26\] CPU.registerFile\[26\]\[26\] _07492_ VGND VGND
+ VPWR VPWR _08193_ sky130_fd_sc_hd__mux2_1
X_10988_ net2149 _05702_ _06190_ VGND VGND VPWR VPWR _06196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18303_ clknet_leaf_12_clk _02583_ VGND VGND VPWR VPWR CPU.PC\[3\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_139_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15515_ _08401_ _03006_ _03009_ _02844_ VGND VGND VPWR VPWR _03010_ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13946__232 clknet_1_0__leaf__07226_ VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__inv_2
X_12727_ _07207_ net1843 _07205_ VGND VGND VPWR VPWR _07208_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_139_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18234_ net75 _02514_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_822 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15446_ _05406_ VGND VGND VPWR VPWR _02943_ sky130_fd_sc_hd__clkbuf_8
X_12658_ net1490 _07154_ VGND VGND VPWR VPWR _00022_ sky130_fd_sc_hd__xor2_1
XFILLER_0_154_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18165_ clknet_leaf_29_clk _02445_ VGND VGND VPWR VPWR CPU.aluIn1\[31\] sky130_fd_sc_hd__dfxtp_2
X_14007__288 clknet_1_1__leaf__08360_ VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__inv_2
X_11609_ net1376 _06494_ _06543_ _06539_ VGND VGND VPWR VPWR _01737_ sky130_fd_sc_hd__o211a_1
X_15377_ _02874_ VGND VGND VPWR VPWR _02875_ sky130_fd_sc_hd__buf_6
XFILLER_0_154_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12589_ net1615 _05425_ _07084_ VGND VGND VPWR VPWR _07118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_10_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_8
X_17116_ clknet_leaf_18_clk _00018_ VGND VGND VPWR VPWR CPU.cycles\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_152_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14200__378 clknet_1_0__leaf__08429_ VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__inv_2
X_18096_ net159 _02376_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[26\] sky130_fd_sc_hd__dfxtp_1
Xhold406 CPU.registerFile\[14\]\[0\] VGND VGND VPWR VPWR net1647 sky130_fd_sc_hd__dlygate4sd3_1
Xhold417 CPU.registerFile\[2\]\[24\] VGND VGND VPWR VPWR net1658 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold428 CPU.registerFile\[11\]\[30\] VGND VGND VPWR VPWR net1669 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold439 CPU.registerFile\[6\]\[23\] VGND VGND VPWR VPWR net1680 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__02705_ clknet_0__02705_ VGND VGND VPWR VPWR clknet_1_1__leaf__02705_
+ sky130_fd_sc_hd__clkbuf_16
X_17047_ net305 _01369_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14259_ _05318_ _05351_ _05367_ _08437_ VGND VGND VPWR VPWR _08438_ sky130_fd_sc_hd__or4b_1
XFILLER_0_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_746 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14354__492 clknet_1_1__leaf__08468_ VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_55_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ CPU.aluIn1\[6\] CPU.Bimm\[6\] VGND VGND VPWR VPWR _04540_ sky130_fd_sc_hd__nor2_1
Xclkbuf_0__02667_ _02667_ VGND VGND VPWR VPWR clknet_0__02667_ sky130_fd_sc_hd__clkbuf_16
X_13992__274 clknet_1_1__leaf__08359_ VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__inv_2
Xhold1106 CPU.registerFile\[15\]\[29\] VGND VGND VPWR VPWR net2347 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1117 CPU.registerFile\[8\]\[11\] VGND VGND VPWR VPWR net2358 sky130_fd_sc_hd__dlygate4sd3_1
X_08751_ _04470_ _04231_ VGND VGND VPWR VPWR _04471_ sky130_fd_sc_hd__nor2_1
Xhold1128 CPU.registerFile\[21\]\[9\] VGND VGND VPWR VPWR net2369 sky130_fd_sc_hd__dlygate4sd3_1
X_17949_ net1138 _02233_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[29\] sky130_fd_sc_hd__dfxtp_1
Xhold1139 CPU.registerFile\[12\]\[7\] VGND VGND VPWR VPWR net2380 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_136_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08682_ _04268_ CPU.aluIn1\[9\] VGND VGND VPWR VPWR _04402_ sky130_fd_sc_hd__and2b_1
XFILLER_0_136_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09303_ _04782_ _05010_ _04777_ VGND VGND VPWR VPWR _05011_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09234_ _04242_ _04944_ VGND VGND VPWR VPWR _04945_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_146_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09165_ CPU.PC\[3\] _04868_ VGND VGND VPWR VPWR _04877_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09096_ _04217_ VGND VGND VPWR VPWR _04808_ sky130_fd_sc_hd__clkbuf_4
X_14437__567 clknet_1_0__leaf__02659_ VGND VGND VPWR VPWR net599 sky130_fd_sc_hd__inv_2
XFILLER_0_102_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold940 CPU.registerFile\[15\]\[2\] VGND VGND VPWR VPWR net2181 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold951 CPU.registerFile\[22\]\[3\] VGND VGND VPWR VPWR net2192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 CPU.registerFile\[6\]\[14\] VGND VGND VPWR VPWR net2203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold973 CPU.registerFile\[20\]\[5\] VGND VGND VPWR VPWR net2214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold984 CPU.registerFile\[31\]\[23\] VGND VGND VPWR VPWR net2225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 CPU.registerFile\[30\]\[5\] VGND VGND VPWR VPWR net2236 sky130_fd_sc_hd__dlygate4sd3_1
X_09998_ _05553_ net1560 _05558_ VGND VGND VPWR VPWR _05592_ sky130_fd_sc_hd__mux2_1
X_08949_ net1706 _04659_ _04668_ VGND VGND VPWR VPWR _04669_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_48_Left_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11960_ _04659_ net1807 _06747_ VGND VGND VPWR VPWR _06748_ sky130_fd_sc_hd__mux2_1
X_14903__987 clknet_1_1__leaf__02705_ VGND VGND VPWR VPWR net1019 sky130_fd_sc_hd__inv_2
X_10911_ _06155_ VGND VGND VPWR VPWR _02051_ sky130_fd_sc_hd__clkbuf_1
X_14602__715 clknet_1_1__leaf__02676_ VGND VGND VPWR VPWR net747 sky130_fd_sc_hd__inv_2
X_11891_ _06710_ VGND VGND VPWR VPWR _06711_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_86_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13630_ CPU.registerFile\[2\]\[22\] _07322_ VGND VGND VPWR VPWR _08051_ sky130_fd_sc_hd__or2_1
X_10842_ _06118_ VGND VGND VPWR VPWR _02083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__02656_ clknet_0__02656_ VGND VGND VPWR VPWR clknet_1_0__leaf__02656_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_39_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13561_ CPU.rs2\[19\] _07705_ _07969_ _07984_ _07737_ VGND VGND VPWR VPWR _01314_
+ sky130_fd_sc_hd__o221a_1
X_10773_ _05511_ net1603 _06081_ VGND VGND VPWR VPWR _06082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_323 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15300_ CPU.registerFile\[27\]\[0\] CPU.registerFile\[31\]\[0\] _02798_ VGND VGND
+ VPWR VPWR _02799_ sky130_fd_sc_hd__mux2_1
X_12512_ _07077_ VGND VGND VPWR VPWR _01334_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16280_ _02818_ _03752_ _03753_ _03227_ VGND VGND VPWR VPWR _03754_ sky130_fd_sc_hd__a22o_1
X_15009__1082 clknet_1_0__leaf__02716_ VGND VGND VPWR VPWR net1114 sky130_fd_sc_hd__inv_2
X_13492_ CPU.registerFile\[5\]\[17\] CPU.registerFile\[4\]\[17\] _04985_ VGND VGND
+ VPWR VPWR _07918_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_57_Left_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12443_ _05306_ net2057 _07035_ VGND VGND VPWR VPWR _07041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_117_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12374_ _07004_ VGND VGND VPWR VPWR _01399_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_134_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14113_ _04660_ _05235_ _00000_ VGND VGND VPWR VPWR _08385_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11325_ _05518_ net2171 _06371_ VGND VGND VPWR VPWR _06375_ sky130_fd_sc_hd__mux2_1
X_15093_ _07185_ _02733_ _02727_ VGND VGND VPWR VPWR _02276_ sky130_fd_sc_hd__a21oi_1
X_15050__1117 clknet_1_0__leaf__02721_ VGND VGND VPWR VPWR net1149 sky130_fd_sc_hd__inv_2
X_11256_ _06338_ VGND VGND VPWR VPWR _01889_ sky130_fd_sc_hd__clkbuf_1
X_10207_ _05714_ VGND VGND VPWR VPWR _02329_ sky130_fd_sc_hd__clkbuf_1
X_11187_ _05516_ net2141 _06299_ VGND VGND VPWR VPWR _06302_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_66_Left_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17803_ net992 _02087_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_10138_ net1732 _05448_ _05632_ VGND VGND VPWR VPWR _05667_ sky130_fd_sc_hd__mux2_1
X_15995_ _02949_ _03473_ _03476_ VGND VGND VPWR VPWR _03477_ sky130_fd_sc_hd__or3_4
X_17734_ net923 _02018_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[20\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_50_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10069_ net2152 _05448_ _05595_ VGND VGND VPWR VPWR _05630_ sky130_fd_sc_hd__mux2_1
X_17665_ net854 _01953_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_14878__964 clknet_1_0__leaf__02703_ VGND VGND VPWR VPWR net996 sky130_fd_sc_hd__inv_2
X_16616_ _03983_ VGND VGND VPWR VPWR _02545_ sky130_fd_sc_hd__clkbuf_1
X_13828_ _07370_ _08242_ VGND VGND VPWR VPWR _08243_ sky130_fd_sc_hd__or2_1
X_17596_ net785 _01884_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13759_ CPU.registerFile\[1\]\[26\] _07576_ _08175_ _07639_ VGND VGND VPWR VPWR _08176_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_75_Left_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16478_ _03195_ _03943_ _03944_ _03945_ _08396_ VGND VGND VPWR VPWR _03946_ sky130_fd_sc_hd__a221o_1
XFILLER_0_155_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18217_ net58 _02497_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15429_ _02760_ VGND VGND VPWR VPWR _02926_ sky130_fd_sc_hd__buf_4
XFILLER_0_26_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18148_ clknet_leaf_19_clk _02428_ VGND VGND VPWR VPWR CPU.aluIn1\[14\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold203 mapped_spi_ram.rcv_data\[2\] VGND VGND VPWR VPWR net1444 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold214 _02183_ VGND VGND VPWR VPWR net1455 sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 per_uart.uart0.enable16_counter\[7\] VGND VGND VPWR VPWR net1466 sky130_fd_sc_hd__dlygate4sd3_1
X_18079_ net142 _02359_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[9\] sky130_fd_sc_hd__dfxtp_1
Xhold236 _02194_ VGND VGND VPWR VPWR net1477 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold247 _07153_ VGND VGND VPWR VPWR net1488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 _00003_ VGND VGND VPWR VPWR net1499 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ _05380_ VGND VGND VPWR VPWR _05549_ sky130_fd_sc_hd__clkbuf_8
Xhold269 CPU.cycles\[28\] VGND VGND VPWR VPWR net1510 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_84_Left_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09852_ _05502_ VGND VGND VPWR VPWR _02504_ sky130_fd_sc_hd__clkbuf_1
X_08803_ CPU.Iimm\[0\] CPU.Bimm\[11\] CPU.instr\[5\] VGND VGND VPWR VPWR _04523_ sky130_fd_sc_hd__mux2_4
XFILLER_0_147_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09783_ net2351 _04958_ _05452_ VGND VGND VPWR VPWR _05462_ sky130_fd_sc_hd__mux2_1
X_08734_ CPU.rs2\[20\] _04201_ _04206_ VGND VGND VPWR VPWR _04454_ sky130_fd_sc_hd__a21oi_1
X_08665_ _04384_ VGND VGND VPWR VPWR _04385_ sky130_fd_sc_hd__inv_2
XANTENNA_109 _05406_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08596_ _04315_ VGND VGND VPWR VPWR _04316_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_93_Left_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09217_ CPU.PC\[22\] CPU.PC\[21\] _04928_ VGND VGND VPWR VPWR _04929_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_622 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09148_ CPU.PC\[8\] CPU.Bimm\[8\] _04820_ VGND VGND VPWR VPWR _04860_ sky130_fd_sc_hd__and3_1
X_14370__507 clknet_1_1__leaf__02652_ VGND VGND VPWR VPWR net539 sky130_fd_sc_hd__inv_2
XFILLER_0_102_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09079_ _04671_ _04788_ _04791_ _04678_ VGND VGND VPWR VPWR _04792_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11110_ CPU.registerFile\[8\]\[23\] _05687_ _06252_ VGND VGND VPWR VPWR _06261_ sky130_fd_sc_hd__mux2_1
X_12090_ _05426_ net2029 _06782_ VGND VGND VPWR VPWR _06816_ sky130_fd_sc_hd__mux2_1
X_15133__1162 clknet_1_0__leaf__02744_ VGND VGND VPWR VPWR net1194 sky130_fd_sc_hd__inv_2
Xhold770 CPU.registerFile\[1\]\[31\] VGND VGND VPWR VPWR net2011 sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 CPU.registerFile\[4\]\[31\] VGND VGND VPWR VPWR net2022 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_112_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11041_ net1660 _05687_ _06215_ VGND VGND VPWR VPWR _06224_ sky130_fd_sc_hd__mux2_1
Xhold792 CPU.registerFile\[25\]\[19\] VGND VGND VPWR VPWR net2033 sky130_fd_sc_hd__dlygate4sd3_1
X_15780_ _02759_ _03265_ _03267_ _02767_ VGND VGND VPWR VPWR _03268_ sky130_fd_sc_hd__a211o_1
X_12992_ CPU.registerFile\[21\]\[3\] _07244_ _07429_ CPU.registerFile\[17\]\[3\] _07431_
+ VGND VGND VPWR VPWR _07432_ sky130_fd_sc_hd__o221a_1
X_11943_ _06738_ VGND VGND VPWR VPWR _01599_ sky130_fd_sc_hd__clkbuf_1
X_17450_ net639 _01738_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14662_ clknet_1_1__leaf__02675_ VGND VGND VPWR VPWR _02682_ sky130_fd_sc_hd__buf_1
X_11874_ net1950 _05721_ _06697_ VGND VGND VPWR VPWR _06702_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__02708_ clknet_0__02708_ VGND VGND VPWR VPWR clknet_1_0__leaf__02708_
+ sky130_fd_sc_hd__clkbuf_16
X_16401_ CPU.registerFile\[20\]\[29\] _02855_ _03026_ VGND VGND VPWR VPWR _03871_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_95_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13613_ CPU.registerFile\[21\]\[21\] _07281_ _07521_ CPU.registerFile\[17\]\[21\]
+ _04972_ VGND VGND VPWR VPWR _08035_ sky130_fd_sc_hd__o221a_1
X_17381_ net570 _01669_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_10825_ _06109_ VGND VGND VPWR VPWR _02091_ sky130_fd_sc_hd__clkbuf_1
X_16332_ CPU.registerFile\[5\]\[27\] CPU.registerFile\[4\]\[27\] _02805_ VGND VGND
+ VPWR VPWR _03804_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_119_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13544_ _07380_ _07963_ _07967_ _07646_ VGND VGND VPWR VPWR _07968_ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10756_ _05495_ net1851 _06070_ VGND VGND VPWR VPWR _06073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16263_ CPU.registerFile\[13\]\[25\] _02889_ _02764_ _03736_ VGND VGND VPWR VPWR
+ _03737_ sky130_fd_sc_hd__o211a_1
X_13475_ CPU.registerFile\[15\]\[17\] _07281_ _07521_ CPU.registerFile\[11\]\[17\]
+ _07253_ VGND VGND VPWR VPWR _07901_ sky130_fd_sc_hd__o221a_1
X_10687_ _06036_ VGND VGND VPWR VPWR _02156_ sky130_fd_sc_hd__clkbuf_1
X_18002_ net1175 _00004_ VGND VGND VPWR VPWR mapped_spi_flash.state\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_152_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12426_ _05130_ net2084 _07024_ VGND VGND VPWR VPWR _07032_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16194_ CPU.registerFile\[6\]\[23\] _03026_ _02763_ _03669_ VGND VGND VPWR VPWR _03670_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12357_ _06995_ VGND VGND VPWR VPWR _01407_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11308_ _05501_ net1940 _06360_ VGND VGND VPWR VPWR _06366_ sky130_fd_sc_hd__mux2_1
X_12288_ _06951_ VGND VGND VPWR VPWR _01432_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_52_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11239_ _06329_ VGND VGND VPWR VPWR _01897_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_147_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15978_ _05010_ _03457_ _03460_ VGND VGND VPWR VPWR _03461_ sky130_fd_sc_hd__or3_2
XFILLER_0_26_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14466__593 clknet_1_0__leaf__02662_ VGND VGND VPWR VPWR net625 sky130_fd_sc_hd__inv_2
X_17717_ net906 _02001_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_14929_ clknet_1_0__leaf__02708_ VGND VGND VPWR VPWR _02709_ sky130_fd_sc_hd__buf_1
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17648_ net837 _01936_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17579_ net768 _01867_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09002_ _04681_ _04718_ _04655_ VGND VGND VPWR VPWR _04719_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_115_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14631__741 clknet_1_1__leaf__02679_ VGND VGND VPWR VPWR net773 sky130_fd_sc_hd__inv_2
XFILLER_0_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09904_ _05537_ net2511 _05533_ VGND VGND VPWR VPWR _05538_ sky130_fd_sc_hd__mux2_1
X_09835_ _05490_ VGND VGND VPWR VPWR _05491_ sky130_fd_sc_hd__buf_4
X_14549__668 clknet_1_1__leaf__02670_ VGND VGND VPWR VPWR net700 sky130_fd_sc_hd__inv_2
X_15008__1081 clknet_1_0__leaf__02716_ VGND VGND VPWR VPWR net1113 sky130_fd_sc_hd__inv_2
X_09766_ _05453_ VGND VGND VPWR VPWR _02541_ sky130_fd_sc_hd__clkbuf_1
X_08717_ _04329_ _04258_ VGND VGND VPWR VPWR _04437_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09697_ _05275_ _05383_ _05387_ _05286_ VGND VGND VPWR VPWR _05388_ sky130_fd_sc_hd__o211a_1
Xrebuffer40 net1282 VGND VGND VPWR VPWR net1281 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_83_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08648_ _04224_ _04365_ _04367_ VGND VGND VPWR VPWR _04368_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_96_658 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08579_ _04196_ _04197_ _04198_ _04298_ VGND VGND VPWR VPWR _04299_ sky130_fd_sc_hd__a211o_1
X_10610_ mapped_spi_flash.rcv_data\[17\] _05981_ VGND VGND VPWR VPWR _05988_ sky130_fd_sc_hd__or2_1
X_11590_ net1372 _06517_ _06509_ _06531_ VGND VGND VPWR VPWR _06532_ sky130_fd_sc_hd__a211o_1
XFILLER_0_25_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10541_ _05940_ VGND VGND VPWR VPWR _02205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14714__816 clknet_1_1__leaf__02687_ VGND VGND VPWR VPWR net848 sky130_fd_sc_hd__inv_2
XFILLER_0_91_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14294__438 clknet_1_0__leaf__08462_ VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__inv_2
X_13260_ CPU.registerFile\[31\]\[10\] _07482_ _07692_ _07621_ _07483_ VGND VGND VPWR
+ VPWR _07693_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_98_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10472_ net1397 _05850_ _05851_ _05883_ VGND VGND VPWR VPWR _05884_ sky130_fd_sc_hd__a211o_1
XFILLER_0_150_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12211_ _06892_ VGND VGND VPWR VPWR _01450_ sky130_fd_sc_hd__clkbuf_1
X_13191_ _07418_ _07624_ _07625_ VGND VGND VPWR VPWR _07626_ sky130_fd_sc_hd__o21a_1
X_12142_ _05230_ net1823 _06841_ VGND VGND VPWR VPWR _06844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16950_ net245 _01276_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_12073_ _06807_ VGND VGND VPWR VPWR _01537_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11024_ _06214_ VGND VGND VPWR VPWR _06215_ sky130_fd_sc_hd__buf_4
X_15901_ CPU.registerFile\[2\]\[14\] _03143_ _02980_ CPU.registerFile\[3\]\[14\] _03144_
+ VGND VGND VPWR VPWR _03386_ sky130_fd_sc_hd__a221o_1
X_16881_ _03973_ _04153_ VGND VGND VPWR VPWR _04164_ sky130_fd_sc_hd__and2b_1
X_15832_ CPU.registerFile\[6\]\[12\] _03057_ _03140_ _03318_ VGND VGND VPWR VPWR _03319_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_129_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14760__858 clknet_1_1__leaf__02691_ VGND VGND VPWR VPWR net890 sky130_fd_sc_hd__inv_2
X_15763_ _05361_ VGND VGND VPWR VPWR _03252_ sky130_fd_sc_hd__buf_4
XFILLER_0_87_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12975_ _07412_ _07413_ _07415_ VGND VGND VPWR VPWR _07416_ sky130_fd_sc_hd__o21a_1
X_16520__188 clknet_1_1__leaf__03963_ VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__inv_2
X_17502_ net691 _01790_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_11926_ _06729_ VGND VGND VPWR VPWR _01607_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_142_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15694_ _02827_ _03183_ _03184_ VGND VGND VPWR VPWR _03185_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_142_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ net622 net1323 VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[26\] sky130_fd_sc_hd__dfxtp_1
X_11857_ CPU.registerFile\[10\]\[15\] _05704_ _06686_ VGND VGND VPWR VPWR _06693_
+ sky130_fd_sc_hd__mux2_1
X_17364_ net553 _01652_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10808_ _05547_ net1859 _06092_ VGND VGND VPWR VPWR _06100_ sky130_fd_sc_hd__mux2_1
X_11788_ _06656_ VGND VGND VPWR VPWR _01672_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16315_ CPU.registerFile\[22\]\[26\] _03032_ VGND VGND VPWR VPWR _03788_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_31_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13527_ _07268_ _07948_ _07951_ VGND VGND VPWR VPWR _07952_ sky130_fd_sc_hd__or3_1
X_17295_ net484 _01583_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_10739_ _06063_ VGND VGND VPWR VPWR _02131_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16246_ _03717_ _03718_ _03720_ _02812_ VGND VGND VPWR VPWR _03721_ sky130_fd_sc_hd__o22a_1
XFILLER_0_153_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13458_ _07474_ _07881_ _07884_ VGND VGND VPWR VPWR _07885_ sky130_fd_sc_hd__or3_1
XFILLER_0_125_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12409_ _04958_ net2301 _07013_ VGND VGND VPWR VPWR _07023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_140_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16177_ CPU.registerFile\[22\]\[22\] CPU.registerFile\[23\]\[22\] _03066_ VGND VGND
+ VPWR VPWR _03654_ sky130_fd_sc_hd__mux2_1
X_13389_ _07272_ VGND VGND VPWR VPWR _07818_ sky130_fd_sc_hd__buf_4
XFILLER_0_23_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_121_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_149_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09620_ _04637_ _05310_ _05313_ _05308_ VGND VGND VPWR VPWR _05314_ sky130_fd_sc_hd__o22a_1
X_09551_ _05245_ _05247_ _04374_ VGND VGND VPWR VPWR _05248_ sky130_fd_sc_hd__mux2_1
X_08502_ CPU.aluIn1\[30\] _04221_ VGND VGND VPWR VPWR _04222_ sky130_fd_sc_hd__nand2_1
XFILLER_0_144_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09482_ _04319_ _04323_ VGND VGND VPWR VPWR _05182_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_65_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16495__165 clknet_1_0__leaf__02756_ VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__inv_2
XFILLER_0_78_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15132__1161 clknet_1_1__leaf__02744_ VGND VGND VPWR VPWR net1193 sky130_fd_sc_hd__inv_2
XFILLER_0_59_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14482__608 clknet_1_0__leaf__02663_ VGND VGND VPWR VPWR net640 sky130_fd_sc_hd__inv_2
X_09818_ _05480_ VGND VGND VPWR VPWR _02516_ sky130_fd_sc_hd__clkbuf_1
X_09749_ _04211_ _05428_ _05430_ _05437_ VGND VGND VPWR VPWR _05438_ sky130_fd_sc_hd__a211o_1
XFILLER_0_68_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_124_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ mapped_spi_ram.rcv_data\[6\] _06601_ VGND VGND VPWR VPWR _06610_ sky130_fd_sc_hd__or2_1
X_12691_ CPU.cycles\[30\] _07172_ VGND VGND VPWR VPWR _07175_ sky130_fd_sc_hd__or2_1
X_11642_ net1521 _06562_ _06567_ VGND VGND VPWR VPWR _01728_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14302__445 clknet_1_1__leaf__08463_ VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__inv_2
XFILLER_0_119_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11573_ _06512_ _05900_ VGND VGND VPWR VPWR _06520_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_30_Left_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16100_ _03252_ _03570_ _03578_ _02935_ VGND VGND VPWR VPWR _03579_ sky130_fd_sc_hd__o211a_1
X_13312_ CPU.registerFile\[21\]\[12\] _07244_ _07429_ CPU.registerFile\[17\]\[12\]
+ _07742_ VGND VGND VPWR VPWR _07743_ sky130_fd_sc_hd__o221a_1
X_10524_ _05926_ _04535_ VGND VGND VPWR VPWR _05928_ sky130_fd_sc_hd__and2b_1
X_17080_ net338 _01402_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_761 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16031_ CPU.registerFile\[29\]\[18\] _02918_ VGND VGND VPWR VPWR _03512_ sky130_fd_sc_hd__or2_1
X_13243_ CPU.registerFile\[6\]\[10\] CPU.registerFile\[7\]\[10\] _07641_ VGND VGND
+ VPWR VPWR _07676_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10455_ CPU.aluIn1\[14\] _04496_ _05868_ VGND VGND VPWR VPWR _05869_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13174_ _07392_ _07604_ _07608_ _07232_ VGND VGND VPWR VPWR _07609_ sky130_fd_sc_hd__o211a_1
X_10386_ _04192_ VGND VGND VPWR VPWR _05816_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12125_ net1244 net2372 _06830_ VGND VGND VPWR VPWR _06835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17982_ net1170 _02266_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_12056_ _06798_ VGND VGND VPWR VPWR _01545_ sky130_fd_sc_hd__clkbuf_1
X_16933_ clknet_leaf_9_clk _01259_ VGND VGND VPWR VPWR per_uart.uart0.txd_reg\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_11007_ net1791 _05721_ _06201_ VGND VGND VPWR VPWR _06206_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_144_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16864_ _04151_ _03976_ _03975_ VGND VGND VPWR VPWR _04152_ sky130_fd_sc_hd__o21ba_1
X_15815_ _02759_ _03299_ _03301_ _02767_ VGND VGND VPWR VPWR _03302_ sky130_fd_sc_hd__a211o_1
X_16795_ _04101_ _04105_ _05815_ VGND VGND VPWR VPWR _02602_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15746_ CPU.registerFile\[20\]\[10\] _02855_ _03026_ VGND VGND VPWR VPWR _03235_
+ sky130_fd_sc_hd__a21o_1
X_12958_ _04937_ VGND VGND VPWR VPWR _07399_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_47_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11909_ _06720_ VGND VGND VPWR VPWR _01615_ sky130_fd_sc_hd__clkbuf_1
X_15677_ CPU.registerFile\[30\]\[8\] CPU.registerFile\[26\]\[8\] _02787_ VGND VGND
+ VPWR VPWR _03168_ sky130_fd_sc_hd__mux2_1
XANTENNA_270 _05509_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12889_ CPU.registerFile\[16\]\[1\] CPU.registerFile\[20\]\[1\] _07314_ VGND VGND
+ VPWR VPWR _07331_ sky130_fd_sc_hd__mux2_1
XANTENNA_281 _05551_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_292 _07232_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17416_ net605 _01704_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14578__694 clknet_1_0__leaf__02673_ VGND VGND VPWR VPWR net726 sky130_fd_sc_hd__inv_2
X_17347_ net536 _01635_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_60_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15007__1080 clknet_1_0__leaf__02716_ VGND VGND VPWR VPWR net1112 sky130_fd_sc_hd__inv_2
X_17278_ net467 _01566_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_796 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16229_ CPU.registerFile\[9\]\[24\] _02802_ _03125_ VGND VGND VPWR VPWR _03704_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_58_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08982_ _04224_ _04698_ _04699_ _04225_ VGND VGND VPWR VPWR _04700_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_143_Right_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14743__842 clknet_1_0__leaf__02690_ VGND VGND VPWR VPWR net874 sky130_fd_sc_hd__inv_2
X_09603_ _04278_ _04312_ VGND VGND VPWR VPWR _05298_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16503__172 clknet_1_0__leaf__03962_ VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__inv_2
Xwire20 _04125_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_1
X_09534_ _05231_ VGND VGND VPWR VPWR _02559_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09465_ _04892_ _05165_ VGND VGND VPWR VPWR _05166_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_708 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_149_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09396_ _04440_ _05099_ VGND VGND VPWR VPWR _05100_ sky130_fd_sc_hd__and2b_1
XFILLER_0_47_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10240_ _05736_ VGND VGND VPWR VPWR _02318_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10171_ net2107 _05689_ _05671_ VGND VGND VPWR VPWR _05690_ sky130_fd_sc_hd__mux2_1
X_14826__917 clknet_1_1__leaf__02698_ VGND VGND VPWR VPWR net949 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_110_Right_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13930_ _07818_ _08340_ _08341_ VGND VGND VPWR VPWR _08342_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_109_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13861_ _07273_ _08273_ _08274_ VGND VGND VPWR VPWR _08275_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_1_0__f__08463_ clknet_0__08463_ VGND VGND VPWR VPWR clknet_1_0__leaf__08463_
+ sky130_fd_sc_hd__clkbuf_16
X_15600_ CPU.registerFile\[28\]\[6\] _02791_ VGND VGND VPWR VPWR _03093_ sky130_fd_sc_hd__or2_1
X_12812_ _05283_ net14 VGND VGND VPWR VPWR _07255_ sky130_fd_sc_hd__nor2_4
XFILLER_0_69_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13792_ _07801_ _08205_ _08206_ _08207_ _07555_ VGND VGND VPWR VPWR _08208_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_122_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15531_ _02819_ VGND VGND VPWR VPWR _03026_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_97_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12743_ _07218_ VGND VGND VPWR VPWR _01262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_139_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_814 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18250_ net91 _02530_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_15462_ _07228_ VGND VGND VPWR VPWR _02958_ sky130_fd_sc_hd__buf_2
X_12674_ CPU.cycles\[22\] _07162_ net1437 VGND VGND VPWR VPWR _07165_ sky130_fd_sc_hd__a21oi_1
X_14872__959 clknet_1_1__leaf__02702_ VGND VGND VPWR VPWR net991 sky130_fd_sc_hd__inv_2
X_17201_ clknet_leaf_11_clk _01489_ VGND VGND VPWR VPWR CPU.Bimm\[12\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18181_ net212 _02461_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[15\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_42_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11625_ mapped_spi_ram.state\[2\] mapped_spi_ram.state\[0\] mapped_spi_ram.state\[1\]
+ _06487_ net2 VGND VGND VPWR VPWR _06555_ sky130_fd_sc_hd__o311a_2
XFILLER_0_5_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_42_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15393_ _02885_ _02886_ _02888_ _02890_ _08396_ VGND VGND VPWR VPWR _02891_ sky130_fd_sc_hd__o221a_1
XFILLER_0_64_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17132_ clknet_leaf_22_clk _00035_ VGND VGND VPWR VPWR CPU.cycles\[28\] sky130_fd_sc_hd__dfxtp_1
X_11556_ net1390 _06499_ _06489_ _06506_ VGND VGND VPWR VPWR _06507_ sky130_fd_sc_hd__a211o_1
XFILLER_0_80_675 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17063_ net321 _01385_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_10507_ net1391 _05892_ _05913_ _05885_ VGND VGND VPWR VPWR _02212_ sky130_fd_sc_hd__o211a_1
Xclkbuf_1_1__f__02721_ clknet_0__02721_ VGND VGND VPWR VPWR clknet_1_1__leaf__02721_
+ sky130_fd_sc_hd__clkbuf_16
X_14275_ _08453_ VGND VGND VPWR VPWR _08454_ sky130_fd_sc_hd__clkbuf_2
X_11487_ _05543_ net2407 _06455_ VGND VGND VPWR VPWR _06461_ sky130_fd_sc_hd__mux2_1
X_16014_ _03491_ _03495_ _02810_ VGND VGND VPWR VPWR _03496_ sky130_fd_sc_hd__a21o_1
X_13226_ CPU.registerFile\[29\]\[9\] _07414_ _07326_ CPU.registerFile\[25\]\[9\] _07489_
+ VGND VGND VPWR VPWR _07660_ sky130_fd_sc_hd__o221a_1
Xclkbuf_0__02752_ _02752_ VGND VGND VPWR VPWR clknet_0__02752_ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_1__f__02652_ clknet_0__02652_ VGND VGND VPWR VPWR clknet_1_1__leaf__02652_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10438_ mapped_spi_flash.cmd_addr\[19\] _04592_ _05820_ VGND VGND VPWR VPWR _05857_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13157_ _07474_ _07589_ _07592_ VGND VGND VPWR VPWR _07593_ sky130_fd_sc_hd__or3_1
Xclkbuf_0__02683_ _02683_ VGND VGND VPWR VPWR clknet_0__02683_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_21_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10369_ _05806_ VGND VGND VPWR VPWR _02244_ sky130_fd_sc_hd__clkbuf_1
X_15131__1160 clknet_1_0__leaf__02744_ VGND VGND VPWR VPWR net1192 sky130_fd_sc_hd__inv_2
X_12108_ _04780_ net1754 _06819_ VGND VGND VPWR VPWR _06826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13088_ CPU.registerFile\[31\]\[5\] _07289_ _07290_ CPU.registerFile\[27\]\[5\] _07345_
+ VGND VGND VPWR VPWR _07526_ sky130_fd_sc_hd__o221a_1
X_17965_ net1153 _02249_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12039_ _06789_ VGND VGND VPWR VPWR _01553_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16916_ net1819 _04182_ VGND VGND VPWR VPWR _04187_ sky130_fd_sc_hd__or2_1
X_17896_ net1085 _02180_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[14\] sky130_fd_sc_hd__dfxtp_1
X_16847_ net2069 net2224 _04139_ VGND VGND VPWR VPWR _04142_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16778_ _04032_ net1763 VGND VGND VPWR VPWR _04091_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15729_ _05093_ _03216_ _03217_ _03218_ _03028_ VGND VGND VPWR VPWR _03219_ sky130_fd_sc_hd__o221a_1
X_09250_ _04385_ _04449_ _04343_ VGND VGND VPWR VPWR _04960_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_118_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_157_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09181_ CPU.PC\[12\] _04851_ VGND VGND VPWR VPWR _04893_ sky130_fd_sc_hd__or2_1
XFILLER_0_146_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_1__f__03968_ clknet_0__03968_ VGND VGND VPWR VPWR clknet_1_1__leaf__03968_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_43_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__08357_ clknet_0__08357_ VGND VGND VPWR VPWR clknet_1_1__leaf__08357_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_73_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08965_ _04222_ _04683_ VGND VGND VPWR VPWR _04684_ sky130_fd_sc_hd__nor2_1
X_14331__471 clknet_1_0__leaf__08466_ VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__inv_2
X_08896_ _04594_ _04599_ VGND VGND VPWR VPWR _04616_ sky130_fd_sc_hd__and2b_1
XFILLER_0_98_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclone3 _05065_ VGND VGND VPWR VPWR net1244 sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_88_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__02672_ clknet_0__02672_ VGND VGND VPWR VPWR clknet_1_0__leaf__02672_
+ sky130_fd_sc_hd__clkbuf_16
X_09517_ _04428_ _04403_ _04427_ VGND VGND VPWR VPWR _05215_ sky130_fd_sc_hd__nor3_1
XFILLER_0_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14594__709 clknet_1_1__leaf__02674_ VGND VGND VPWR VPWR net741 sky130_fd_sc_hd__inv_2
XFILLER_0_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09448_ _05149_ VGND VGND VPWR VPWR _05150_ sky130_fd_sc_hd__buf_4
XFILLER_0_94_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_149_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09379_ _04843_ _04900_ VGND VGND VPWR VPWR _05084_ sky130_fd_sc_hd__and2b_1
XFILLER_0_46_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11410_ _06420_ VGND VGND VPWR VPWR _01817_ sky130_fd_sc_hd__clkbuf_1
X_12390_ _07012_ VGND VGND VPWR VPWR _07013_ sky130_fd_sc_hd__buf_4
XFILLER_0_62_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11341_ _06383_ VGND VGND VPWR VPWR _01849_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12772__221 clknet_1_0__leaf__07225_ VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_104_Left_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11272_ CPU.registerFile\[9\]\[11\] _05712_ _06346_ VGND VGND VPWR VPWR _06347_ sky130_fd_sc_hd__mux2_1
X_14414__546 clknet_1_0__leaf__02657_ VGND VGND VPWR VPWR net578 sky130_fd_sc_hd__inv_2
XFILLER_0_30_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13011_ CPU.registerFile\[28\]\[3\] CPU.registerFile\[24\]\[3\] _07297_ VGND VGND
+ VPWR VPWR _07451_ sky130_fd_sc_hd__mux2_1
X_10223_ _05332_ VGND VGND VPWR VPWR _05725_ sky130_fd_sc_hd__clkbuf_4
X_10154_ _05678_ VGND VGND VPWR VPWR _02346_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17750_ net939 _02034_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_14962_ clknet_1_0__leaf__02708_ VGND VGND VPWR VPWR _02712_ sky130_fd_sc_hd__buf_1
X_10085_ _05639_ VGND VGND VPWR VPWR _02376_ sky130_fd_sc_hd__clkbuf_1
X_16701_ _03991_ net2289 VGND VGND VPWR VPWR _04026_ sky130_fd_sc_hd__nand2_1
Xclkbuf_1_0__f__03988_ clknet_0__03988_ VGND VGND VPWR VPWR clknet_1_0__leaf__03988_
+ sky130_fd_sc_hd__clkbuf_16
X_13913_ CPU.registerFile\[6\]\[31\] CPU.registerFile\[7\]\[31\] _07641_ VGND VGND
+ VPWR VPWR _08325_ sky130_fd_sc_hd__mux2_1
X_17681_ net870 _01969_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[3\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_113_Left_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13844_ CPU.registerFile\[6\]\[28\] CPU.registerFile\[7\]\[28\] _07311_ VGND VGND
+ VPWR VPWR _08259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13775_ _07412_ _08190_ _08191_ VGND VGND VPWR VPWR _08192_ sky130_fd_sc_hd__o21a_1
X_10987_ _06195_ VGND VGND VPWR VPWR _02015_ sky130_fd_sc_hd__clkbuf_1
X_18302_ clknet_leaf_12_clk _02582_ VGND VGND VPWR VPWR CPU.PC\[2\] sky130_fd_sc_hd__dfxtp_2
X_14460__588 clknet_1_1__leaf__02661_ VGND VGND VPWR VPWR net620 sky130_fd_sc_hd__inv_2
X_15514_ _08405_ _03007_ _03008_ VGND VGND VPWR VPWR _03009_ sky130_fd_sc_hd__a21o_1
XFILLER_0_84_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12726_ per_uart.d_in_uart\[5\] _07178_ _07203_ per_uart.uart0.txd_reg\[6\] VGND
+ VGND VPWR VPWR _07207_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16494_ net2476 _07228_ _03942_ _03961_ _06482_ VGND VGND VPWR VPWR _02445_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_139_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15445_ CPU.registerFile\[5\]\[2\] CPU.registerFile\[4\]\[2\] _02805_ VGND VGND VPWR
+ VPWR _02942_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_139_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18233_ net74 _02513_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12657_ _07154_ _07155_ VGND VGND VPWR VPWR _00021_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_834 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11608_ net1362 _06501_ _06496_ CPU.mem_wdata\[4\] _06508_ VGND VGND VPWR VPWR _06543_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_142_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18164_ clknet_leaf_29_clk _02444_ VGND VGND VPWR VPWR CPU.aluIn1\[30\] sky130_fd_sc_hd__dfxtp_2
X_15376_ _02854_ VGND VGND VPWR VPWR _02874_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_143_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12588_ _07117_ VGND VGND VPWR VPWR _01265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_122_Left_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17115_ clknet_leaf_18_clk _00017_ VGND VGND VPWR VPWR CPU.cycles\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_152_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18095_ net158 _02375_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_11539_ net1393 _06491_ _06494_ net1326 _05844_ VGND VGND VPWR VPWR _01758_ sky130_fd_sc_hd__o221a_1
XFILLER_0_20_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold407 CPU.registerFile\[14\]\[2\] VGND VGND VPWR VPWR net1648 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold418 CPU.registerFile\[30\]\[30\] VGND VGND VPWR VPWR net1659 sky130_fd_sc_hd__dlygate4sd3_1
X_17046_ net304 _01368_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_150_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14258_ _04411_ _04300_ _05417_ _05428_ _05395_ VGND VGND VPWR VPWR _08437_ sky130_fd_sc_hd__a221oi_1
Xhold429 CPU.registerFile\[28\]\[14\] VGND VGND VPWR VPWR net1670 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__02704_ clknet_0__02704_ VGND VGND VPWR VPWR clknet_1_1__leaf__02704_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13209_ CPU.registerFile\[2\]\[9\] _07322_ VGND VGND VPWR VPWR _07643_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14389__523 clknet_1_1__leaf__02655_ VGND VGND VPWR VPWR net555 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_55_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__02666_ _02666_ VGND VGND VPWR VPWR clknet_0__02666_ sky130_fd_sc_hd__clkbuf_16
X_08750_ CPU.aluIn1\[26\] VGND VGND VPWR VPWR _04470_ sky130_fd_sc_hd__inv_2
Xhold1107 CPU.registerFile\[13\]\[5\] VGND VGND VPWR VPWR net2348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1118 CPU.registerFile\[7\]\[12\] VGND VGND VPWR VPWR net2359 sky130_fd_sc_hd__dlygate4sd3_1
X_17948_ net1137 _02232_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[28\] sky130_fd_sc_hd__dfxtp_1
Xhold1129 CPU.registerFile\[2\]\[19\] VGND VGND VPWR VPWR net2370 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_131_Left_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08681_ _04263_ CPU.aluIn1\[10\] VGND VGND VPWR VPWR _04401_ sky130_fd_sc_hd__and2b_1
XFILLER_0_136_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17879_ net1068 _02163_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_bitcount\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09302_ mapped_spi_ram.rcv_data\[11\] _04783_ _04784_ mapped_spi_flash.rcv_data\[11\]
+ VGND VGND VPWR VPWR _05010_ sky130_fd_sc_hd__a22oi_4
X_14855__943 clknet_1_0__leaf__02701_ VGND VGND VPWR VPWR net975 sky130_fd_sc_hd__inv_2
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09233_ _04244_ _04346_ VGND VGND VPWR VPWR _04944_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09164_ _04873_ _04875_ VGND VGND VPWR VPWR _04876_ sky130_fd_sc_hd__or2b_1
XFILLER_0_17_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09095_ _04461_ _04806_ VGND VGND VPWR VPWR _04807_ sky130_fd_sc_hd__nor2_1
Xhold930 CPU.registerFile\[23\]\[18\] VGND VGND VPWR VPWR net2171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 CPU.registerFile\[3\]\[30\] VGND VGND VPWR VPWR net2182 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold952 CPU.registerFile\[12\]\[27\] VGND VGND VPWR VPWR net2193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold963 CPU.registerFile\[13\]\[22\] VGND VGND VPWR VPWR net2204 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold974 CPU.registerFile\[21\]\[24\] VGND VGND VPWR VPWR net2215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 CPU.registerFile\[27\]\[8\] VGND VGND VPWR VPWR net2226 sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 CPU.registerFile\[22\]\[5\] VGND VGND VPWR VPWR net2237 sky130_fd_sc_hd__dlygate4sd3_1
X_09997_ _05591_ VGND VGND VPWR VPWR _02448_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_4_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08948_ _04667_ VGND VGND VPWR VPWR _04668_ sky130_fd_sc_hd__buf_4
XFILLER_0_99_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08879_ _04590_ _04596_ _04597_ _04598_ CPU.PC\[22\] VGND VGND VPWR VPWR _04599_
+ sky130_fd_sc_hd__a32o_2
X_10910_ net1564 _05691_ _06154_ VGND VGND VPWR VPWR _06155_ sky130_fd_sc_hd__mux2_1
X_11890_ _05450_ _06250_ VGND VGND VPWR VPWR _06710_ sky130_fd_sc_hd__nor2_2
Xclkbuf_1_0__f__02724_ clknet_0__02724_ VGND VGND VPWR VPWR clknet_1_0__leaf__02724_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_157_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10841_ net1822 _05691_ _06117_ VGND VGND VPWR VPWR _06118_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__02655_ clknet_0__02655_ VGND VGND VPWR VPWR clknet_1_0__leaf__02655_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13560_ _07306_ _07976_ _07983_ _07703_ VGND VGND VPWR VPWR _07984_ sky130_fd_sc_hd__a31o_1
Xsplit34 CPU.instr\[5\] VGND VGND VPWR VPWR net1275 sky130_fd_sc_hd__buf_6
X_10772_ _06069_ VGND VGND VPWR VPWR _06081_ sky130_fd_sc_hd__buf_4
X_12511_ net1867 _05723_ _07071_ VGND VGND VPWR VPWR _07077_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13491_ _07915_ _07916_ _07315_ VGND VGND VPWR VPWR _07917_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15230_ clknet_1_0__leaf__02749_ VGND VGND VPWR VPWR _02754_ sky130_fd_sc_hd__buf_1
X_12442_ _07040_ VGND VGND VPWR VPWR _01367_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12373_ _05273_ net1893 _06999_ VGND VGND VPWR VPWR _07004_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14112_ _04647_ _00000_ _08384_ VGND VGND VPWR VPWR _01465_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11324_ _06374_ VGND VGND VPWR VPWR _01857_ sky130_fd_sc_hd__clkbuf_1
X_15092_ net1352 _07184_ VGND VGND VPWR VPWR _02733_ sky130_fd_sc_hd__nand2_1
X_14043_ clknet_1_1__leaf__08363_ VGND VGND VPWR VPWR _08365_ sky130_fd_sc_hd__buf_1
X_11255_ CPU.registerFile\[9\]\[19\] _05696_ _06335_ VGND VGND VPWR VPWR _06338_ sky130_fd_sc_hd__mux2_1
X_10206_ net1967 _05712_ _05713_ VGND VGND VPWR VPWR _05714_ sky130_fd_sc_hd__mux2_1
X_11186_ _06301_ VGND VGND VPWR VPWR _01922_ sky130_fd_sc_hd__clkbuf_1
X_17802_ net991 _02086_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_10137_ _05666_ VGND VGND VPWR VPWR _02351_ sky130_fd_sc_hd__clkbuf_1
X_15994_ _02901_ _03474_ _03475_ _02867_ VGND VGND VPWR VPWR _03476_ sky130_fd_sc_hd__a22o_1
X_15239__148 clknet_1_0__leaf__02754_ VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__inv_2
X_17733_ net922 _02017_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[19\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_50_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10068_ _05629_ VGND VGND VPWR VPWR _02383_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_50_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17664_ net853 _01952_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_14013__293 clknet_1_1__leaf__08361_ VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__inv_2
X_16615_ net1565 net1552 _03979_ VGND VGND VPWR VPWR _03983_ sky130_fd_sc_hd__mux2_1
X_13827_ CPU.registerFile\[28\]\[28\] CPU.registerFile\[24\]\[28\] _04936_ VGND VGND
+ VPWR VPWR _08242_ sky130_fd_sc_hd__mux2_1
X_17595_ net784 _01883_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[13\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_0__f__08429_ clknet_0__08429_ VGND VGND VPWR VPWR clknet_1_0__leaf__08429_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_57_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13758_ CPU.registerFile\[5\]\[26\] CPU.registerFile\[4\]\[26\] _07262_ VGND VGND
+ VPWR VPWR _08175_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12709_ net1351 _07190_ VGND VGND VPWR VPWR _07191_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16477_ CPU.registerFile\[10\]\[31\] _02928_ _02910_ VGND VGND VPWR VPWR _03945_
+ sky130_fd_sc_hd__o21a_1
X_13689_ _07272_ _08108_ VGND VGND VPWR VPWR _08109_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18216_ net57 _02496_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15428_ CPU.registerFile\[27\]\[2\] CPU.registerFile\[31\]\[2\] _02852_ VGND VGND
+ VPWR VPWR _02925_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14994__1069 clknet_1_1__leaf__02714_ VGND VGND VPWR VPWR net1101 sky130_fd_sc_hd__inv_2
XFILLER_0_122_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15359_ _02850_ _02853_ _02856_ VGND VGND VPWR VPWR _02857_ sky130_fd_sc_hd__mux2_1
X_18147_ clknet_leaf_19_clk _02427_ VGND VGND VPWR VPWR CPU.aluIn1\[13\] sky130_fd_sc_hd__dfxtp_4
XFILLER_0_25_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold204 per_uart.uart0.enable16_counter\[11\] VGND VGND VPWR VPWR net1445 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold215 mapped_spi_ram.rcv_data\[4\] VGND VGND VPWR VPWR net1456 sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 CPU.cycles\[3\] VGND VGND VPWR VPWR net1467 sky130_fd_sc_hd__dlygate4sd3_1
X_18078_ net141 _02358_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold237 mapped_spi_ram.rcv_data\[20\] VGND VGND VPWR VPWR net1478 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09920_ _05548_ VGND VGND VPWR VPWR _02482_ sky130_fd_sc_hd__clkbuf_1
Xhold248 CPU.cycles\[27\] VGND VGND VPWR VPWR net1489 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17029_ net287 _01351_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[23\] sky130_fd_sc_hd__dfxtp_1
Xhold259 mapped_spi_flash.rcv_data\[2\] VGND VGND VPWR VPWR net1500 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__02718_ _02718_ VGND VGND VPWR VPWR clknet_0__02718_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09851_ _05501_ net2310 _05491_ VGND VGND VPWR VPWR _05502_ sky130_fd_sc_hd__mux2_1
X_08802_ CPU.aluIn1\[3\] _04521_ VGND VGND VPWR VPWR _04522_ sky130_fd_sc_hd__or2_4
X_09782_ _05461_ VGND VGND VPWR VPWR _02533_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08733_ CPU.aluIn1\[21\] VGND VGND VPWR VPWR _04453_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08664_ _04383_ _04247_ VGND VGND VPWR VPWR _04384_ sky130_fd_sc_hd__nor2_1
XFILLER_0_68_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_68_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08595_ CPU.aluIn1\[8\] _04270_ VGND VGND VPWR VPWR _04315_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_101_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14443__572 clknet_1_1__leaf__02660_ VGND VGND VPWR VPWR net604 sky130_fd_sc_hd__inv_2
X_14181__360 clknet_1_1__leaf__08428_ VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__inv_2
XFILLER_0_9_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09216_ CPU.PC\[20\] _04927_ VGND VGND VPWR VPWR _04928_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_686 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09147_ CPU.PC\[9\] _04858_ VGND VGND VPWR VPWR _04859_ sky130_fd_sc_hd__xor2_1
XFILLER_0_16_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09078_ _04351_ _04790_ _04671_ VGND VGND VPWR VPWR _04791_ sky130_fd_sc_hd__o21ai_1
Xhold760 CPU.registerFile\[30\]\[22\] VGND VGND VPWR VPWR net2001 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_875 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold771 CPU.registerFile\[31\]\[1\] VGND VGND VPWR VPWR net2012 sky130_fd_sc_hd__dlygate4sd3_1
Xhold782 CPU.registerFile\[8\]\[16\] VGND VGND VPWR VPWR net2023 sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ _06223_ VGND VGND VPWR VPWR _01990_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_112_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold793 CPU.registerFile\[19\]\[17\] VGND VGND VPWR VPWR net2034 sky130_fd_sc_hd__dlygate4sd3_1
X_12991_ _07245_ _07430_ VGND VGND VPWR VPWR _07431_ sky130_fd_sc_hd__or2_1
X_14526__647 clknet_1_0__leaf__02668_ VGND VGND VPWR VPWR net679 sky130_fd_sc_hd__inv_2
X_11942_ net2197 _05721_ _06733_ VGND VGND VPWR VPWR _06738_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11873_ _06701_ VGND VGND VPWR VPWR _01632_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__02707_ clknet_0__02707_ VGND VGND VPWR VPWR clknet_1_0__leaf__02707_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13612_ CPU.registerFile\[16\]\[21\] CPU.registerFile\[20\]\[21\] _07785_ VGND VGND
+ VPWR VPWR _08034_ sky130_fd_sc_hd__mux2_1
X_16400_ CPU.registerFile\[22\]\[29\] _08399_ VGND VGND VPWR VPWR _03870_ sky130_fd_sc_hd__and2_1
X_10824_ net1674 _05675_ _06106_ VGND VGND VPWR VPWR _06109_ sky130_fd_sc_hd__mux2_1
X_17380_ net569 _01668_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13543_ _07369_ _07964_ _07966_ _07570_ VGND VGND VPWR VPWR _07967_ sky130_fd_sc_hd__a211o_1
X_16331_ _03195_ _03800_ _03802_ _02965_ VGND VGND VPWR VPWR _03803_ sky130_fd_sc_hd__a211o_1
XFILLER_0_55_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10755_ _06072_ VGND VGND VPWR VPWR _02124_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16262_ CPU.registerFile\[9\]\[25\] _02777_ VGND VGND VPWR VPWR _03736_ sky130_fd_sc_hd__or2_1
X_13474_ CPU.registerFile\[14\]\[17\] CPU.registerFile\[10\]\[17\] _07274_ VGND VGND
+ VPWR VPWR _07900_ sky130_fd_sc_hd__mux2_1
X_10686_ _05493_ net1662 _06034_ VGND VGND VPWR VPWR _06036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18001_ clknet_leaf_7_clk _02285_ VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[15\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12425_ _07031_ VGND VGND VPWR VPWR _01375_ sky130_fd_sc_hd__clkbuf_1
X_16193_ CPU.registerFile\[7\]\[23\] _03317_ VGND VGND VPWR VPWR _03669_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14572__689 clknet_1_0__leaf__02672_ VGND VGND VPWR VPWR net721 sky130_fd_sc_hd__inv_2
X_12356_ _05109_ net1908 _06988_ VGND VGND VPWR VPWR _06995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11307_ _06365_ VGND VGND VPWR VPWR _01865_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15075_ clknet_1_1__leaf__02720_ VGND VGND VPWR VPWR _02724_ sky130_fd_sc_hd__buf_1
X_12287_ CPU.aluReg\[8\] _06950_ _06924_ VGND VGND VPWR VPWR _06951_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_52_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11238_ net1944 _05679_ _06324_ VGND VGND VPWR VPWR _06329_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11169_ _06292_ VGND VGND VPWR VPWR _01930_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_147_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_147_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15977_ _02926_ _03458_ _03459_ VGND VGND VPWR VPWR _03460_ sky130_fd_sc_hd__o21a_1
XFILLER_0_89_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17716_ net905 _02000_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14928_ clknet_1_1__leaf__07222_ VGND VGND VPWR VPWR _02708_ sky130_fd_sc_hd__buf_1
XFILLER_0_117_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17647_ net836 _01935_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17578_ net767 _01866_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09001_ mapped_spi_ram.rcv_data\[4\] _04689_ _04691_ mapped_spi_flash.rcv_data\[4\]
+ VGND VGND VPWR VPWR _04718_ sky130_fd_sc_hd__a22o_2
XFILLER_0_6_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09903_ _05229_ VGND VGND VPWR VPWR _05537_ sky130_fd_sc_hd__buf_4
XFILLER_0_6_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09834_ _05488_ _05489_ VGND VGND VPWR VPWR _05490_ sky130_fd_sc_hd__nand2_4
X_09765_ net2128 _04659_ _05452_ VGND VGND VPWR VPWR _05453_ sky130_fd_sc_hd__mux2_1
X_08716_ _04398_ _04434_ _04435_ VGND VGND VPWR VPWR _04436_ sky130_fd_sc_hd__o21a_1
X_09696_ _05384_ _05281_ _05386_ _05277_ VGND VGND VPWR VPWR _05387_ sky130_fd_sc_hd__o22a_1
Xrebuffer30 net1279 VGND VGND VPWR VPWR net1271 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_68_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer41 net1283 VGND VGND VPWR VPWR net1282 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_83_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08647_ _04222_ _04366_ VGND VGND VPWR VPWR _04367_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_83_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08578_ CPU.mem_wdata\[1\] VGND VGND VPWR VPWR _04298_ sky130_fd_sc_hd__inv_2
XFILLER_0_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10540_ _05830_ _05939_ VGND VGND VPWR VPWR _05940_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_33_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10471_ _05852_ _05882_ VGND VGND VPWR VPWR _05883_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_157_Right_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_134_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12210_ net2514 _06890_ _06891_ VGND VGND VPWR VPWR _06892_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13190_ CPU.registerFile\[13\]\[8\] _07482_ _07420_ CPU.registerFile\[9\]\[8\] _07249_
+ VGND VGND VPWR VPWR _07625_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_131_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12141_ _06843_ VGND VGND VPWR VPWR _01505_ sky130_fd_sc_hd__clkbuf_1
X_12072_ _05209_ CPU.registerFile\[26\]\[10\] _06805_ VGND VGND VPWR VPWR _06807_
+ sky130_fd_sc_hd__mux2_1
Xhold590 CPU.registerFile\[14\]\[27\] VGND VGND VPWR VPWR net1831 sky130_fd_sc_hd__dlygate4sd3_1
X_11023_ _05450_ _06141_ VGND VGND VPWR VPWR _06214_ sky130_fd_sc_hd__nor2_4
X_15900_ CPU.registerFile\[6\]\[14\] _03057_ _03140_ _03384_ VGND VGND VPWR VPWR _03385_
+ sky130_fd_sc_hd__o211a_1
X_16880_ _04163_ VGND VGND VPWR VPWR _02629_ sky130_fd_sc_hd__clkbuf_1
X_15831_ CPU.registerFile\[7\]\[12\] _03317_ VGND VGND VPWR VPWR _03318_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_129_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14993__1068 clknet_1_1__leaf__02714_ VGND VGND VPWR VPWR net1100 sky130_fd_sc_hd__inv_2
X_12974_ CPU.registerFile\[15\]\[2\] _07414_ _07326_ CPU.registerFile\[11\]\[2\] _07252_
+ VGND VGND VPWR VPWR _07415_ sky130_fd_sc_hd__o221a_1
X_15762_ _02924_ _03248_ _03249_ _03250_ _02930_ VGND VGND VPWR VPWR _03251_ sky130_fd_sc_hd__a221o_1
Xhold1290 CPU.registerFile\[15\]\[6\] VGND VGND VPWR VPWR net2531 sky130_fd_sc_hd__dlygate4sd3_1
X_17501_ net690 _01789_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_11925_ CPU.registerFile\[11\]\[15\] _05704_ _06722_ VGND VGND VPWR VPWR _06729_
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_142_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15693_ CPU.registerFile\[18\]\[8\] _02833_ _02836_ CPU.registerFile\[19\]\[8\] _02758_
+ VGND VGND VPWR VPWR _03184_ sky130_fd_sc_hd__o221a_1
XFILLER_0_157_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17432_ net621 _01720_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[25\] sky130_fd_sc_hd__dfxtp_1
X_16579__51 clknet_1_1__leaf__03969_ VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__inv_2
X_11856_ _06692_ VGND VGND VPWR VPWR _01640_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10807_ _06099_ VGND VGND VPWR VPWR _02099_ sky130_fd_sc_hd__clkbuf_1
X_17363_ net552 _01651_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_11787_ _05090_ net1955 _06650_ VGND VGND VPWR VPWR _06656_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_901 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16594__65 clknet_1_1__leaf__03970_ VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__inv_2
X_16314_ CPU.registerFile\[21\]\[26\] CPU.registerFile\[23\]\[26\] _02769_ VGND VGND
+ VPWR VPWR _03787_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13526_ _07475_ _07949_ _07950_ VGND VGND VPWR VPWR _07951_ sky130_fd_sc_hd__o21a_1
X_10738_ _05545_ net2130 _06056_ VGND VGND VPWR VPWR _06063_ sky130_fd_sc_hd__mux2_1
X_17294_ net483 _01582_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16245_ CPU.registerFile\[1\]\[24\] _02939_ _03719_ _02894_ VGND VGND VPWR VPWR _03720_
+ sky130_fd_sc_hd__a22o_1
X_13457_ CPU.registerFile\[27\]\[16\] _07363_ _07883_ VGND VGND VPWR VPWR _07884_
+ sky130_fd_sc_hd__o21a_1
X_10669_ _05964_ _06024_ VGND VGND VPWR VPWR _06025_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_124_Right_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12408_ _07022_ VGND VGND VPWR VPWR _01383_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13388_ _07646_ _07806_ _07809_ _07816_ VGND VGND VPWR VPWR _07817_ sky130_fd_sc_hd__a31o_1
X_16176_ CPU.registerFile\[16\]\[22\] _02833_ _02836_ CPU.registerFile\[17\]\[22\]
+ _02856_ VGND VGND VPWR VPWR _03653_ sky130_fd_sc_hd__o221a_1
XFILLER_0_23_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12339_ _04933_ net2079 _06977_ VGND VGND VPWR VPWR _06986_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_149_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14009_ clknet_1_0__leaf__07223_ VGND VGND VPWR VPWR _08361_ sky130_fd_sc_hd__buf_1
XFILLER_0_37_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14509__631 clknet_1_1__leaf__02667_ VGND VGND VPWR VPWR net663 sky130_fd_sc_hd__inv_2
XFILLER_0_128_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09550_ _04427_ _05246_ VGND VGND VPWR VPWR _05247_ sky130_fd_sc_hd__nor2_1
X_08501_ CPU.rs2\[30\] _04201_ _04206_ VGND VGND VPWR VPWR _04221_ sky130_fd_sc_hd__a21o_1
X_09481_ _04321_ _04214_ _04681_ CPU.aluReg\[11\] _05180_ VGND VGND VPWR VPWR _05181_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_19_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_898 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14555__673 clknet_1_1__leaf__02671_ VGND VGND VPWR VPWR net705 sky130_fd_sc_hd__inv_2
XFILLER_0_132_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09817_ net2279 _05306_ _05474_ VGND VGND VPWR VPWR _05480_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09748_ _05434_ _05436_ _04483_ VGND VGND VPWR VPWR _05437_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14720__821 clknet_1_0__leaf__02688_ VGND VGND VPWR VPWR net853 sky130_fd_sc_hd__inv_2
X_09679_ _04672_ _05367_ _05370_ _04768_ VGND VGND VPWR VPWR _05371_ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11710_ net1481 _06603_ _06609_ _06607_ VGND VGND VPWR VPWR _01702_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_124_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12690_ CPU.cycles\[30\] _07172_ VGND VGND VPWR VPWR _07174_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11641_ _06499_ _06555_ _06566_ VGND VGND VPWR VPWR _06567_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14638__748 clknet_1_0__leaf__02679_ VGND VGND VPWR VPWR net780 sky130_fd_sc_hd__inv_2
X_11572_ net1358 _06495_ _06519_ _06516_ VGND VGND VPWR VPWR _01750_ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13311_ _07245_ _07741_ VGND VGND VPWR VPWR _07742_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10523_ _04518_ _04634_ _05926_ _04629_ VGND VGND VPWR VPWR _05927_ sky130_fd_sc_hd__a31o_1
XFILLER_0_91_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13242_ CPU.registerFile\[1\]\[10\] _07576_ _07674_ _07639_ VGND VGND VPWR VPWR _07675_
+ sky130_fd_sc_hd__a22o_1
X_16030_ CPU.registerFile\[27\]\[18\] CPU.registerFile\[31\]\[18\] _03050_ VGND VGND
+ VPWR VPWR _03511_ sky130_fd_sc_hd__mux2_1
X_10454_ _04553_ _04556_ _04555_ VGND VGND VPWR VPWR _05868_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13173_ _07288_ _07607_ VGND VGND VPWR VPWR _07608_ sky130_fd_sc_hd__or2_1
X_10385_ _05812_ net1329 _05813_ net2539 _05815_ VGND VGND VPWR VPWR _02237_ sky130_fd_sc_hd__a221o_1
X_12124_ _06834_ VGND VGND VPWR VPWR _01513_ sky130_fd_sc_hd__clkbuf_1
X_17981_ net1169 _02265_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12055_ net1245 net1785 _06794_ VGND VGND VPWR VPWR _06798_ sky130_fd_sc_hd__mux2_1
X_16932_ clknet_leaf_9_clk _01258_ VGND VGND VPWR VPWR per_uart.uart0.txd_reg\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_11006_ _06205_ VGND VGND VPWR VPWR _02006_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_144_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16863_ per_uart.uart0.uart_rxd2 VGND VGND VPWR VPWR _04151_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_144_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14383__518 clknet_1_1__leaf__02654_ VGND VGND VPWR VPWR net550 sky130_fd_sc_hd__inv_2
X_15814_ CPU.registerFile\[8\]\[12\] _02763_ _03117_ _03300_ VGND VGND VPWR VPWR _03301_
+ sky130_fd_sc_hd__o211a_1
X_14949__1028 clknet_1_0__leaf__02710_ VGND VGND VPWR VPWR net1060 sky130_fd_sc_hd__inv_2
X_16794_ _04050_ _04102_ _04103_ _04104_ VGND VGND VPWR VPWR _04105_ sky130_fd_sc_hd__a31o_1
XFILLER_0_88_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15745_ CPU.registerFile\[22\]\[10\] _08399_ VGND VGND VPWR VPWR _03234_ sky130_fd_sc_hd__and2_1
X_12957_ _05338_ VGND VGND VPWR VPWR _07398_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_47_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11908_ CPU.registerFile\[11\]\[23\] _05687_ _06711_ VGND VGND VPWR VPWR _06720_
+ sky130_fd_sc_hd__mux2_1
X_15676_ _03162_ _03166_ _02784_ VGND VGND VPWR VPWR _03167_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12888_ _07291_ VGND VGND VPWR VPWR _07330_ sky130_fd_sc_hd__buf_4
XANTENNA_260 _05050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_271 _05524_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_282 _05551_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17415_ net604 _01703_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[8\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_293 _07268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11839_ _06683_ VGND VGND VPWR VPWR _01648_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17346_ net535 _01634_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_60_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13509_ CPU.registerFile\[2\]\[18\] _07388_ VGND VGND VPWR VPWR _07934_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17277_ net466 _01565_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_155_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_879 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_130_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16228_ CPU.registerFile\[13\]\[24\] _03123_ VGND VGND VPWR VPWR _03703_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_469 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16159_ CPU.registerFile\[15\]\[22\] _02889_ VGND VGND VPWR VPWR _03636_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08981_ _04210_ VGND VGND VPWR VPWR _04699_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_58_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09602_ _04423_ _05296_ VGND VGND VPWR VPWR _05297_ sky130_fd_sc_hd__nor2_1
X_09533_ net2020 _05230_ _05189_ VGND VGND VPWR VPWR _05231_ sky130_fd_sc_hd__mux2_1
X_09464_ _04852_ _04893_ VGND VGND VPWR VPWR _05165_ sky130_fd_sc_hd__and2b_1
XFILLER_0_47_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09395_ _04439_ _04394_ _04438_ VGND VGND VPWR VPWR _05099_ sky130_fd_sc_hd__or3_1
X_16558__32 clknet_1_0__leaf__03967_ VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__inv_2
XFILLER_0_149_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16573__46 clknet_1_0__leaf__03968_ VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__inv_2
XFILLER_0_144_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_879 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14992__1067 clknet_1_1__leaf__02714_ VGND VGND VPWR VPWR net1099 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_95_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10170_ _04957_ VGND VGND VPWR VPWR _05689_ sky130_fd_sc_hd__buf_2
XFILLER_0_30_776 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14219__395 clknet_1_0__leaf__08431_ VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__inv_2
XFILLER_0_100_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13860_ CPU.registerFile\[23\]\[29\] _07361_ _07283_ CPU.registerFile\[19\]\[29\]
+ _07253_ VGND VGND VPWR VPWR _08274_ sky130_fd_sc_hd__o221a_1
Xclkbuf_1_0__f__08462_ clknet_0__08462_ VGND VGND VPWR VPWR clknet_1_0__leaf__08462_
+ sky130_fd_sc_hd__clkbuf_16
X_12811_ _07253_ VGND VGND VPWR VPWR _07254_ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_2_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13791_ CPU.registerFile\[3\]\[27\] _07804_ _07987_ VGND VGND VPWR VPWR _08207_ sky130_fd_sc_hd__o21a_1
X_15530_ _02854_ VGND VGND VPWR VPWR _03025_ sky130_fd_sc_hd__buf_4
X_12742_ _07217_ net1698 _07205_ VGND VGND VPWR VPWR _07218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12673_ CPU.cycles\[22\] CPU.cycles\[23\] _07162_ VGND VGND VPWR VPWR _07164_ sky130_fd_sc_hd__and3_1
X_15461_ CPU.aluIn1\[2\] _07705_ _02933_ _02957_ _07737_ VGND VGND VPWR VPWR _02416_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_155_826 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_843 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17200_ clknet_leaf_11_clk _01488_ VGND VGND VPWR VPWR CPU.Bimm\[10\] sky130_fd_sc_hd__dfxtp_4
X_11624_ _06493_ _06552_ _06553_ _06470_ VGND VGND VPWR VPWR _06554_ sky130_fd_sc_hd__a31o_1
X_18180_ net211 _02460_ VGND VGND VPWR VPWR CPU.registerFile\[14\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_42_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15392_ CPU.registerFile\[27\]\[1\] _02889_ _02780_ VGND VGND VPWR VPWR _02890_ sky130_fd_sc_hd__a21o_1
XFILLER_0_154_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17131_ clknet_leaf_22_clk _00034_ VGND VGND VPWR VPWR CPU.cycles\[27\] sky130_fd_sc_hd__dfxtp_1
X_11555_ _06501_ _05877_ VGND VGND VPWR VPWR _06506_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10506_ net1382 _05887_ _05856_ _05912_ VGND VGND VPWR VPWR _05913_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_21_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14274_ _08448_ _08449_ _08451_ _08452_ VGND VGND VPWR VPWR _08453_ sky130_fd_sc_hd__a31o_2
X_17062_ net320 _01384_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[24\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__02720_ clknet_0__02720_ VGND VGND VPWR VPWR clknet_1_1__leaf__02720_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_80_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11486_ _06460_ VGND VGND VPWR VPWR _01781_ sky130_fd_sc_hd__clkbuf_1
X_16013_ _02914_ _03492_ _03494_ _02864_ VGND VGND VPWR VPWR _03495_ sky130_fd_sc_hd__a211o_1
X_13225_ CPU.registerFile\[28\]\[9\] CPU.registerFile\[24\]\[9\] _07476_ VGND VGND
+ VPWR VPWR _07659_ sky130_fd_sc_hd__mux2_1
Xclkbuf_0__02751_ _02751_ VGND VGND VPWR VPWR clknet_0__02751_ sky130_fd_sc_hd__clkbuf_16
X_10437_ _05826_ VGND VGND VPWR VPWR _05856_ sky130_fd_sc_hd__buf_2
XFILLER_0_20_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13156_ _07418_ _07590_ _07591_ VGND VGND VPWR VPWR _07592_ sky130_fd_sc_hd__o21a_1
Xclkbuf_0__02682_ _02682_ VGND VGND VPWR VPWR clknet_0__02682_ sky130_fd_sc_hd__clkbuf_16
X_10368_ _05545_ net2362 _05799_ VGND VGND VPWR VPWR _05806_ sky130_fd_sc_hd__mux2_1
X_12107_ _06825_ VGND VGND VPWR VPWR _01521_ sky130_fd_sc_hd__clkbuf_1
X_13087_ _07351_ _07524_ VGND VGND VPWR VPWR _07525_ sky130_fd_sc_hd__or2_1
X_17964_ net1152 _02248_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[9\] sky130_fd_sc_hd__dfxtp_1
X_10299_ _05545_ net2214 _05762_ VGND VGND VPWR VPWR _05769_ sky130_fd_sc_hd__mux2_1
X_12038_ _04762_ net1924 _06783_ VGND VGND VPWR VPWR _06789_ sky130_fd_sc_hd__mux2_1
X_16915_ CPU.mem_wdata\[3\] _04180_ _04186_ _04176_ VGND VGND VPWR VPWR _02641_ sky130_fd_sc_hd__o211a_1
X_17895_ net1084 _02179_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16846_ net1541 VGND VGND VPWR VPWR _02617_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_0_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_743 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16777_ _04086_ _04090_ _05815_ VGND VGND VPWR VPWR _02599_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15728_ CPU.registerFile\[20\]\[9\] _03025_ _03026_ VGND VGND VPWR VPWR _03218_ sky130_fd_sc_hd__a21o_1
X_15659_ CPU.registerFile\[16\]\[7\] _03068_ _03069_ CPU.registerFile\[17\]\[7\] _02779_
+ VGND VGND VPWR VPWR _03151_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_157_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09180_ _04856_ _04891_ _04854_ VGND VGND VPWR VPWR _04892_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17329_ net518 _01617_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[25\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__03967_ clknet_0__03967_ VGND VGND VPWR VPWR clknet_1_1__leaf__03967_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_126_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__08356_ clknet_0__08356_ VGND VGND VPWR VPWR clknet_1_1__leaf__08356_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08964_ _04682_ VGND VGND VPWR VPWR _04683_ sky130_fd_sc_hd__clkbuf_4
X_14667__774 clknet_1_1__leaf__02682_ VGND VGND VPWR VPWR net806 sky130_fd_sc_hd__inv_2
X_08895_ _04601_ _04604_ VGND VGND VPWR VPWR _04615_ sky130_fd_sc_hd__and2_1
Xclone4 _05045_ VGND VGND VPWR VPWR net1245 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f__02671_ clknet_0__02671_ VGND VGND VPWR VPWR clknet_1_0__leaf__02671_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09516_ _04216_ _05212_ _05213_ _05134_ _04717_ VGND VGND VPWR VPWR _05214_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_104_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09447_ _05135_ _05140_ _05148_ VGND VGND VPWR VPWR _05149_ sky130_fd_sc_hd__or3b_4
XFILLER_0_148_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09378_ _05074_ _05075_ _05082_ _04773_ VGND VGND VPWR VPWR _05083_ sky130_fd_sc_hd__o31a_1
X_14832__922 clknet_1_1__leaf__02699_ VGND VGND VPWR VPWR net954 sky130_fd_sc_hd__inv_2
XFILLER_0_47_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11340_ _05532_ net2413 _06382_ VGND VGND VPWR VPWR _06383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14948__1027 clknet_1_0__leaf__02710_ VGND VGND VPWR VPWR net1059 sky130_fd_sc_hd__inv_2
XFILLER_0_132_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11271_ _06323_ VGND VGND VPWR VPWR _06346_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_104_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13010_ CPU.registerFile\[31\]\[3\] _07289_ _07290_ CPU.registerFile\[27\]\[3\] _07449_
+ VGND VGND VPWR VPWR _07450_ sky130_fd_sc_hd__o221a_1
X_10222_ _05724_ VGND VGND VPWR VPWR _02324_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10153_ net1958 _05677_ _05671_ VGND VGND VPWR VPWR _05678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10084_ net2041 _04762_ _05633_ VGND VGND VPWR VPWR _05639_ sky130_fd_sc_hd__mux2_1
X_16700_ _04021_ _04025_ _04015_ VGND VGND VPWR VPWR _02587_ sky130_fd_sc_hd__a21oi_1
X_13912_ net1493 _08018_ _08324_ _08017_ VGND VGND VPWR VPWR _01325_ sky130_fd_sc_hd__o211a_1
X_17680_ net869 _01968_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_13843_ CPU.registerFile\[1\]\[28\] _07256_ _08257_ _07368_ VGND VGND VPWR VPWR _08258_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10986_ net2297 _05700_ _06190_ VGND VGND VPWR VPWR _06195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13774_ CPU.registerFile\[29\]\[26\] _07414_ _07326_ CPU.registerFile\[25\]\[26\]
+ _07489_ VGND VGND VPWR VPWR _08191_ sky130_fd_sc_hd__o221a_1
XFILLER_0_58_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18301_ net35 _02581_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[31\] sky130_fd_sc_hd__dfxtp_1
X_15513_ CPU.registerFile\[2\]\[4\] _02872_ _02873_ CPU.registerFile\[3\]\[4\] _02875_
+ VGND VGND VPWR VPWR _03008_ sky130_fd_sc_hd__a221o_1
X_12725_ _07206_ VGND VGND VPWR VPWR _01256_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_26_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16493_ _02757_ _03951_ _03960_ _07308_ VGND VGND VPWR VPWR _03961_ sky130_fd_sc_hd__a31o_1
XFILLER_0_155_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14495__619 clknet_1_1__leaf__02665_ VGND VGND VPWR VPWR net651 sky130_fd_sc_hd__inv_2
XFILLER_0_127_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_139_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18232_ net73 _02512_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_15444_ CPU.registerFile\[2\]\[2\] _02872_ _02939_ CPU.registerFile\[3\]\[2\] _02940_
+ VGND VGND VPWR VPWR _02941_ sky130_fd_sc_hd__a221o_1
X_16537__13 clknet_1_1__leaf__03965_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__inv_2
X_12656_ net1524 _07152_ VGND VGND VPWR VPWR _07155_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18163_ clknet_leaf_29_clk _02443_ VGND VGND VPWR VPWR CPU.aluIn1\[29\] sky130_fd_sc_hd__dfxtp_2
X_11607_ net1388 _06524_ _06542_ _06539_ VGND VGND VPWR VPWR _01738_ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12587_ net1602 _05401_ _07107_ VGND VGND VPWR VPWR _07117_ sky130_fd_sc_hd__mux2_1
X_15375_ _02822_ VGND VGND VPWR VPWR _02873_ sky130_fd_sc_hd__buf_4
XFILLER_0_5_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17114_ clknet_leaf_18_clk _00016_ VGND VGND VPWR VPWR CPU.cycles\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16552__27 clknet_1_1__leaf__03966_ VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__inv_2
X_18094_ net157 _02374_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_11538_ mapped_spi_ram.state\[2\] _06493_ _06487_ VGND VGND VPWR VPWR _06494_ sky130_fd_sc_hd__o21a_2
XFILLER_0_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold408 CPU.registerFile\[5\]\[25\] VGND VGND VPWR VPWR net1649 sky130_fd_sc_hd__dlygate4sd3_1
Xhold419 CPU.registerFile\[7\]\[23\] VGND VGND VPWR VPWR net1660 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__02703_ clknet_0__02703_ VGND VGND VPWR VPWR clknet_1_1__leaf__02703_
+ sky130_fd_sc_hd__clkbuf_16
X_17045_ net303 _01367_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_11469_ _06451_ VGND VGND VPWR VPWR _01789_ sky130_fd_sc_hd__clkbuf_1
X_14257_ _05288_ VGND VGND VPWR VPWR _08436_ sky130_fd_sc_hd__buf_2
XFILLER_0_151_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13208_ CPU.registerFile\[6\]\[9\] CPU.registerFile\[7\]\[9\] _07641_ VGND VGND VPWR
+ VPWR _07642_ sky130_fd_sc_hd__mux2_1
X_14809__902 clknet_1_1__leaf__02696_ VGND VGND VPWR VPWR net934 sky130_fd_sc_hd__inv_2
XFILLER_0_21_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13139_ _07254_ _07569_ _07574_ _07232_ VGND VGND VPWR VPWR _07575_ sky130_fd_sc_hd__o211a_1
Xclkbuf_0__02665_ _02665_ VGND VGND VPWR VPWR clknet_0__02665_ sky130_fd_sc_hd__clkbuf_16
X_12749__202 clknet_1_0__leaf__07221_ VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__inv_2
Xhold1108 CPU.registerFile\[4\]\[14\] VGND VGND VPWR VPWR net2349 sky130_fd_sc_hd__dlygate4sd3_1
X_17947_ net1136 _02231_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[27\] sky130_fd_sc_hd__dfxtp_1
Xhold1119 CPU.registerFile\[8\]\[24\] VGND VGND VPWR VPWR net2360 sky130_fd_sc_hd__dlygate4sd3_1
X_08680_ _04399_ _04320_ VGND VGND VPWR VPWR _04400_ sky130_fd_sc_hd__nor2_1
X_17878_ net1067 _02162_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_bitcount\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16829_ per_uart.uart0.tx_bitcount\[0\] _04129_ per_uart.uart0.tx_bitcount\[1\] VGND
+ VGND VPWR VPWR _04130_ sky130_fd_sc_hd__mux2_1
X_14991__1066 clknet_1_1__leaf__02714_ VGND VGND VPWR VPWR net1098 sky130_fd_sc_hd__inv_2
X_15216__127 clknet_1_1__leaf__02752_ VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__inv_2
XFILLER_0_88_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09301_ _05009_ VGND VGND VPWR VPWR _02570_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_152_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09232_ _04240_ _04214_ _04808_ CPU.aluReg\[22\] _04942_ VGND VGND VPWR VPWR _04943_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09163_ _04871_ _04874_ VGND VGND VPWR VPWR _04875_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09094_ _04701_ VGND VGND VPWR VPWR _04806_ sky130_fd_sc_hd__buf_2
XFILLER_0_32_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold920 CPU.registerFile\[31\]\[26\] VGND VGND VPWR VPWR net2161 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold931 CPU.registerFile\[30\]\[17\] VGND VGND VPWR VPWR net2172 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold942 CPU.registerFile\[22\]\[11\] VGND VGND VPWR VPWR net2183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold953 CPU.registerFile\[25\]\[26\] VGND VGND VPWR VPWR net2194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold964 CPU.registerFile\[23\]\[1\] VGND VGND VPWR VPWR net2205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold975 CPU.registerFile\[19\]\[27\] VGND VGND VPWR VPWR net2216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold986 CPU.registerFile\[3\]\[14\] VGND VGND VPWR VPWR net2227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold997 CPU.registerFile\[21\]\[29\] VGND VGND VPWR VPWR net2238 sky130_fd_sc_hd__dlygate4sd3_1
X_09996_ _05551_ net1648 _05581_ VGND VGND VPWR VPWR _05591_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_4_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08947_ _04662_ _04666_ VGND VGND VPWR VPWR _04667_ sky130_fd_sc_hd__nor2_4
X_08878_ _04586_ VGND VGND VPWR VPWR _04598_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_0__f__02723_ clknet_0__02723_ VGND VGND VPWR VPWR clknet_1_0__leaf__02723_
+ sky130_fd_sc_hd__clkbuf_16
X_10840_ _06105_ VGND VGND VPWR VPWR _06117_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_1_0__f__02654_ clknet_0__02654_ VGND VGND VPWR VPWR clknet_1_0__leaf__02654_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10771_ _06080_ VGND VGND VPWR VPWR _02116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12510_ _07076_ VGND VGND VPWR VPWR _01335_ sky130_fd_sc_hd__clkbuf_1
X_13490_ CPU.registerFile\[6\]\[17\] CPU.registerFile\[7\]\[17\] _07311_ VGND VGND
+ VPWR VPWR _07916_ sky130_fd_sc_hd__mux2_1
X_14420__551 clknet_1_0__leaf__02658_ VGND VGND VPWR VPWR net583 sky130_fd_sc_hd__inv_2
XFILLER_0_54_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12441_ _05273_ net1877 _07035_ VGND VGND VPWR VPWR _07040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12372_ _07003_ VGND VGND VPWR VPWR _01400_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_782 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14111_ _04661_ _00000_ VGND VGND VPWR VPWR _08384_ sky130_fd_sc_hd__nor2_1
X_11323_ _05516_ net2253 _06371_ VGND VGND VPWR VPWR _06374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15091_ _07184_ _02732_ _02727_ VGND VGND VPWR VPWR _02275_ sky130_fd_sc_hd__a21oi_1
X_14338__478 clknet_1_1__leaf__08466_ VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__inv_2
X_11254_ _06337_ VGND VGND VPWR VPWR _01890_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10205_ _05670_ VGND VGND VPWR VPWR _05713_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_770 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11185_ _05514_ net1729 _06299_ VGND VGND VPWR VPWR _06301_ sky130_fd_sc_hd__mux2_1
X_17801_ net990 _02085_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_10136_ net2085 _05426_ _05632_ VGND VGND VPWR VPWR _05666_ sky130_fd_sc_hd__mux2_1
X_15993_ CPU.registerFile\[19\]\[17\] CPU.registerFile\[17\]\[17\] _03025_ VGND VGND
+ VPWR VPWR _03475_ sky130_fd_sc_hd__mux2_1
X_17732_ net921 _02016_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_10067_ net1963 _05426_ _05595_ VGND VGND VPWR VPWR _05629_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_2_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17663_ net852 _01951_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_14804__898 clknet_1_1__leaf__02695_ VGND VGND VPWR VPWR net930 sky130_fd_sc_hd__inv_2
XFILLER_0_89_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16614_ _03982_ VGND VGND VPWR VPWR _02544_ sky130_fd_sc_hd__clkbuf_1
X_13826_ _08237_ _08240_ _07405_ VGND VGND VPWR VPWR _08241_ sky130_fd_sc_hd__mux2_1
X_17594_ net783 _01882_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_14048__324 clknet_1_0__leaf__08365_ VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__inv_2
X_14503__626 clknet_1_1__leaf__02666_ VGND VGND VPWR VPWR net658 sky130_fd_sc_hd__inv_2
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__08428_ clknet_0__08428_ VGND VGND VPWR VPWR clknet_1_0__leaf__08428_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13757_ CPU.rs2\[25\] _07705_ _08158_ _08174_ _07737_ VGND VGND VPWR VPWR _01320_
+ sky130_fd_sc_hd__o221a_1
X_10969_ net2328 _05683_ _06179_ VGND VGND VPWR VPWR _06186_ sky130_fd_sc_hd__mux2_1
X_14241__414 clknet_1_1__leaf__08434_ VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f__08359_ clknet_0__08359_ VGND VGND VPWR VPWR clknet_1_0__leaf__08359_
+ sky130_fd_sc_hd__clkbuf_16
X_12779__228 clknet_1_0__leaf__07225_ VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__inv_2
X_12708_ net1445 _07189_ VGND VGND VPWR VPWR _07190_ sky130_fd_sc_hd__or2_1
X_16476_ CPU.registerFile\[14\]\[31\] _03072_ VGND VGND VPWR VPWR _03944_ sky130_fd_sc_hd__or2_1
X_13688_ CPU.registerFile\[8\]\[23\] CPU.registerFile\[12\]\[23\] _07265_ VGND VGND
+ VPWR VPWR _08108_ sky130_fd_sc_hd__mux2_1
X_18215_ net56 _02495_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15427_ _02923_ VGND VGND VPWR VPWR _02924_ sky130_fd_sc_hd__buf_4
XFILLER_0_127_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12639_ CPU.cycles\[7\] _07142_ net1496 VGND VGND VPWR VPWR _07145_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18146_ clknet_leaf_19_clk _02426_ VGND VGND VPWR VPWR CPU.aluIn1\[12\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15358_ _02855_ VGND VGND VPWR VPWR _02856_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold205 _02738_ VGND VGND VPWR VPWR net1446 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18077_ net140 _02357_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[7\] sky130_fd_sc_hd__dfxtp_1
Xhold216 per_uart.uart0.enable16_counter\[10\] VGND VGND VPWR VPWR net1457 sky130_fd_sc_hd__dlygate4sd3_1
X_15289_ CPU.registerFile\[30\]\[0\] CPU.registerFile\[26\]\[0\] _02787_ VGND VGND
+ VPWR VPWR _02788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold227 mapped_spi_flash.rcv_data\[26\] VGND VGND VPWR VPWR net1468 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 CPU.rs2\[31\] VGND VGND VPWR VPWR net1479 sky130_fd_sc_hd__dlygate4sd3_1
X_17028_ net286 _01350_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[22\] sky130_fd_sc_hd__dfxtp_1
Xhold249 CPU.cycles\[16\] VGND VGND VPWR VPWR net1490 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_0__02717_ _02717_ VGND VGND VPWR VPWR clknet_0__02717_ sky130_fd_sc_hd__clkbuf_16
X_09850_ _04761_ VGND VGND VPWR VPWR _05501_ sky130_fd_sc_hd__clkbuf_4
X_08801_ CPU.Iimm\[3\] CPU.Bimm\[3\] _04372_ VGND VGND VPWR VPWR _04521_ sky130_fd_sc_hd__mux2_4
X_09781_ net1809 _04933_ _05452_ VGND VGND VPWR VPWR _05461_ sky130_fd_sc_hd__mux2_1
X_08732_ _04449_ _04385_ _04343_ _04451_ VGND VGND VPWR VPWR _04452_ sky130_fd_sc_hd__a211o_1
X_08663_ CPU.aluIn1\[19\] VGND VGND VPWR VPWR _04383_ sky130_fd_sc_hd__inv_2
X_14947__1026 clknet_1_1__leaf__02710_ VGND VGND VPWR VPWR net1058 sky130_fd_sc_hd__inv_2
XFILLER_0_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08594_ _04312_ _04278_ _04313_ _04275_ VGND VGND VPWR VPWR _04314_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_68_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14779__875 clknet_1_1__leaf__02693_ VGND VGND VPWR VPWR net907 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_85_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_138_Right_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09215_ CPU.PC\[19\] CPU.PC\[18\] _04926_ VGND VGND VPWR VPWR _04927_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09146_ CPU.Bimm\[9\] _04820_ VGND VGND VPWR VPWR _04858_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_698 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09077_ _04350_ _04789_ VGND VGND VPWR VPWR _04790_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_116_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold750 CPU.registerFile\[11\]\[24\] VGND VGND VPWR VPWR net1991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold761 CPU.registerFile\[12\]\[24\] VGND VGND VPWR VPWR net2002 sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 CPU.registerFile\[6\]\[11\] VGND VGND VPWR VPWR net2013 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_887 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold783 CPU.registerFile\[19\]\[1\] VGND VGND VPWR VPWR net2024 sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 mapped_spi_flash.rcv_data\[3\] VGND VGND VPWR VPWR net2035 sky130_fd_sc_hd__dlygate4sd3_1
X_09979_ _05582_ VGND VGND VPWR VPWR _02457_ sky130_fd_sc_hd__clkbuf_1
X_12990_ CPU.registerFile\[16\]\[3\] CPU.registerFile\[20\]\[3\] _07240_ VGND VGND
+ VPWR VPWR _07430_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11941_ _06737_ VGND VGND VPWR VPWR _01600_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_28_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ net2367 _05719_ _06697_ VGND VGND VPWR VPWR _06701_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__02706_ clknet_0__02706_ VGND VGND VPWR VPWR clknet_1_0__leaf__02706_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13611_ _08025_ _08032_ _07334_ VGND VGND VPWR VPWR _08033_ sky130_fd_sc_hd__mux2_1
X_10823_ _06108_ VGND VGND VPWR VPWR _02092_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_105_Right_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16330_ CPU.registerFile\[15\]\[27\] _02889_ _02770_ _03801_ VGND VGND VPWR VPWR
+ _03802_ sky130_fd_sc_hd__o211a_1
X_13542_ CPU.registerFile\[3\]\[19\] _07373_ _07965_ _07376_ VGND VGND VPWR VPWR _07966_
+ sky130_fd_sc_hd__o211a_1
X_10754_ _05493_ net1659 _06070_ VGND VGND VPWR VPWR _06072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16261_ CPU.registerFile\[15\]\[25\] CPU.registerFile\[11\]\[25\] _02761_ VGND VGND
+ VPWR VPWR _03735_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13473_ _07653_ _07897_ _07898_ VGND VGND VPWR VPWR _07899_ sky130_fd_sc_hd__o21a_1
X_10685_ _06035_ VGND VGND VPWR VPWR _02157_ sky130_fd_sc_hd__clkbuf_1
X_18000_ clknet_leaf_7_clk _02284_ VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[14\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12424_ _05109_ net2288 _07024_ VGND VGND VPWR VPWR _07031_ sky130_fd_sc_hd__mux2_1
X_16192_ CPU.registerFile\[2\]\[23\] _02821_ _02822_ CPU.registerFile\[3\]\[23\] _02855_
+ VGND VGND VPWR VPWR _03668_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12355_ _06994_ VGND VGND VPWR VPWR _01408_ sky130_fd_sc_hd__clkbuf_1
X_15245__153 clknet_1_1__leaf__02755_ VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__inv_2
X_14990__1065 clknet_1_1__leaf__02714_ VGND VGND VPWR VPWR net1097 sky130_fd_sc_hd__inv_2
XFILLER_0_23_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11306_ _05499_ net1992 _06360_ VGND VGND VPWR VPWR _06365_ sky130_fd_sc_hd__mux2_1
X_12286_ CPU.aluIn1\[8\] _06949_ _06927_ VGND VGND VPWR VPWR _06950_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11237_ _06328_ VGND VGND VPWR VPWR _01898_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_52_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11168_ _05497_ net2309 _06288_ VGND VGND VPWR VPWR _06292_ sky130_fd_sc_hd__mux2_1
X_10119_ _05657_ VGND VGND VPWR VPWR _02360_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_147_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11099_ _06255_ VGND VGND VPWR VPWR _01963_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15976_ CPU.registerFile\[18\]\[16\] _03068_ _03069_ CPU.registerFile\[19\]\[16\]
+ _03074_ VGND VGND VPWR VPWR _03459_ sky130_fd_sc_hd__o221a_1
X_17715_ net904 _01999_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17646_ net835 _01934_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_13809_ CPU.registerFile\[13\]\[27\] _07282_ _08224_ VGND VGND VPWR VPWR _08225_
+ sky130_fd_sc_hd__o21a_1
X_17577_ net766 _01865_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16459_ net2491 _07228_ _03911_ _03927_ _06482_ VGND VGND VPWR VPWR _02444_ sky130_fd_sc_hd__o221a_1
XFILLER_0_73_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09000_ _04716_ _04652_ _04654_ VGND VGND VPWR VPWR _04717_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_91_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18129_ net192 _02409_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[27\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13959__244 clknet_1_1__leaf__08356_ VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__inv_2
XFILLER_0_158_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09902_ _05536_ VGND VGND VPWR VPWR _02488_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09833_ _04665_ _04663_ _04664_ CPU.writeBack VGND VGND VPWR VPWR _05489_ sky130_fd_sc_hd__and4b_2
XFILLER_0_67_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09764_ _05451_ VGND VGND VPWR VPWR _05452_ sky130_fd_sc_hd__buf_4
X_08715_ _04327_ _04260_ VGND VGND VPWR VPWR _04435_ sky130_fd_sc_hd__or2b_1
XFILLER_0_69_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09695_ mapped_spi_flash.rcv_data\[26\] _04784_ _05385_ VGND VGND VPWR VPWR _05386_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_83_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer20 net1262 VGND VGND VPWR VPWR net1261 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer31 _04526_ VGND VGND VPWR VPWR net1272 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer42 net1284 VGND VGND VPWR VPWR net1283 sky130_fd_sc_hd__buf_2
X_08646_ CPU.aluIn1\[30\] _04221_ VGND VGND VPWR VPWR _04366_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_83_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08577_ _04293_ _04294_ net24 _04291_ _04296_ VGND VGND VPWR VPWR _04297_ sky130_fd_sc_hd__a221o_2
XFILLER_0_147_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_833 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10470_ CPU.PC\[13\] _05867_ _05880_ _05881_ VGND VGND VPWR VPWR _05882_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_150_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09129_ _04839_ _04840_ VGND VGND VPWR VPWR _04841_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_131_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12140_ _05209_ net1993 _06841_ VGND VGND VPWR VPWR _06843_ sky130_fd_sc_hd__mux2_1
X_14077__350 clknet_1_0__leaf__08368_ VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__inv_2
XFILLER_0_103_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14532__652 clknet_1_1__leaf__02669_ VGND VGND VPWR VPWR net684 sky130_fd_sc_hd__inv_2
X_12071_ _06806_ VGND VGND VPWR VPWR _01538_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold580 CPU.registerFile\[1\]\[24\] VGND VGND VPWR VPWR net1821 sky130_fd_sc_hd__dlygate4sd3_1
Xhold591 CPU.registerFile\[15\]\[11\] VGND VGND VPWR VPWR net1832 sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ _06213_ VGND VGND VPWR VPWR _01998_ sky130_fd_sc_hd__clkbuf_1
X_15830_ net15 VGND VGND VPWR VPWR _03317_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_129_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15761_ CPU.registerFile\[13\]\[10\] _02775_ VGND VGND VPWR VPWR _03250_ sky130_fd_sc_hd__or2_1
X_14188__367 clknet_1_0__leaf__08428_ VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__inv_2
X_12973_ _07234_ VGND VGND VPWR VPWR _07414_ sky130_fd_sc_hd__clkbuf_8
Xhold1280 CPU.registerFile\[10\]\[4\] VGND VGND VPWR VPWR net2521 sky130_fd_sc_hd__dlygate4sd3_1
X_17500_ net689 _01788_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[14\] sky130_fd_sc_hd__dfxtp_1
Xhold1291 CPU.registerFile\[25\]\[15\] VGND VGND VPWR VPWR net2532 sky130_fd_sc_hd__dlygate4sd3_1
X_11924_ _06728_ VGND VGND VPWR VPWR _01608_ sky130_fd_sc_hd__clkbuf_1
X_15692_ CPU.registerFile\[22\]\[8\] CPU.registerFile\[23\]\[8\] _02829_ VGND VGND
+ VPWR VPWR _03183_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_142_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17431_ net620 _01719_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11855_ net2250 _05702_ _06686_ VGND VGND VPWR VPWR _06692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_362 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_157_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17362_ net551 _01650_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[26\] sky130_fd_sc_hd__dfxtp_1
X_10806_ _05545_ net2236 _06092_ VGND VGND VPWR VPWR _06099_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11786_ _06655_ VGND VGND VPWR VPWR _01673_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16313_ _02848_ _03781_ _03785_ _02843_ VGND VGND VPWR VPWR _03786_ sky130_fd_sc_hd__a211o_1
XFILLER_0_126_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13525_ CPU.registerFile\[29\]\[18\] _07325_ _07500_ CPU.registerFile\[25\]\[18\]
+ _07249_ VGND VGND VPWR VPWR _07950_ sky130_fd_sc_hd__o221a_1
X_17293_ net482 _01581_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_10737_ _06062_ VGND VGND VPWR VPWR _02132_ sky130_fd_sc_hd__clkbuf_1
X_14916__999 clknet_1_0__leaf__02706_ VGND VGND VPWR VPWR net1031 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_11_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16244_ CPU.registerFile\[5\]\[24\] CPU.registerFile\[4\]\[24\] _03146_ VGND VGND
+ VPWR VPWR _03719_ sky130_fd_sc_hd__mux2_1
X_13456_ CPU.registerFile\[31\]\[16\] _07482_ _07882_ _07621_ _07483_ VGND VGND VPWR
+ VPWR _07883_ sky130_fd_sc_hd__o221a_1
X_14615__727 clknet_1_1__leaf__02677_ VGND VGND VPWR VPWR net759 sky130_fd_sc_hd__inv_2
X_10668_ net1346 _05963_ VGND VGND VPWR VPWR _06024_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12407_ _04933_ net2225 _07013_ VGND VGND VPWR VPWR _07022_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16175_ _05050_ _03651_ VGND VGND VPWR VPWR _03652_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10599_ mapped_spi_flash.rcv_data\[22\] _05981_ VGND VGND VPWR VPWR _05982_ sky130_fd_sc_hd__or2_1
X_13387_ _07812_ _07815_ _07514_ VGND VGND VPWR VPWR _07816_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_23_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14946__1025 clknet_1_1__leaf__02710_ VGND VGND VPWR VPWR net1057 sky130_fd_sc_hd__inv_2
X_12338_ _06985_ VGND VGND VPWR VPWR _01416_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_149_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12269_ CPU.aluIn1\[12\] _06936_ _06927_ VGND VGND VPWR VPWR _06937_ sky130_fd_sc_hd__mux2_1
X_15959_ CPU.registerFile\[24\]\[16\] _03130_ _02780_ _03441_ VGND VGND VPWR VPWR
+ _03442_ sky130_fd_sc_hd__o211a_1
X_14661__769 clknet_1_1__leaf__02681_ VGND VGND VPWR VPWR net801 sky130_fd_sc_hd__inv_2
X_08500_ CPU.aluIn1\[31\] _04207_ _04214_ _04219_ CPU.aluReg\[31\] VGND VGND VPWR
+ VPWR _04220_ sky130_fd_sc_hd__a32o_1
X_09480_ _04322_ _04740_ VGND VGND VPWR VPWR _05180_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_19_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17629_ net818 _01917_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_924 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09816_ _05479_ VGND VGND VPWR VPWR _02517_ sky130_fd_sc_hd__clkbuf_1
X_09747_ _04216_ _04208_ _05435_ VGND VGND VPWR VPWR _05436_ sky130_fd_sc_hd__or3_1
X_09678_ _04800_ _05369_ VGND VGND VPWR VPWR _05370_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_38_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ CPU.aluIn1\[24\] _04235_ VGND VGND VPWR VPWR _04349_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_124_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11640_ mapped_spi_ram.snd_bitcount\[1\] mapped_spi_ram.snd_bitcount\[0\] VGND VGND
+ VPWR VPWR _06566_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11571_ net1361 _06517_ _06509_ _06518_ VGND VGND VPWR VPWR _06519_ sky130_fd_sc_hd__a211o_1
XFILLER_0_9_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13310_ CPU.registerFile\[16\]\[12\] CPU.registerFile\[20\]\[12\] _07240_ VGND VGND
+ VPWR VPWR _07741_ sky130_fd_sc_hd__mux2_1
X_10522_ _04537_ _04536_ VGND VGND VPWR VPWR _05926_ sky130_fd_sc_hd__or2b_1
XFILLER_0_18_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13241_ CPU.registerFile\[5\]\[10\] CPU.registerFile\[4\]\[10\] _07262_ VGND VGND
+ VPWR VPWR _07674_ sky130_fd_sc_hd__mux2_1
X_10453_ _04598_ VGND VGND VPWR VPWR _05867_ sky130_fd_sc_hd__buf_2
XFILLER_0_150_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10384_ _05812_ net1329 _05813_ _05814_ _05815_ VGND VGND VPWR VPWR _02238_ sky130_fd_sc_hd__a221oi_1
X_13172_ CPU.registerFile\[21\]\[8\] _07502_ _07503_ CPU.registerFile\[17\]\[8\] _07606_
+ VGND VGND VPWR VPWR _07607_ sky130_fd_sc_hd__o221a_1
XFILLER_0_60_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12123_ net1245 net1854 _06830_ VGND VGND VPWR VPWR _06834_ sky130_fd_sc_hd__mux2_1
X_17980_ net1168 _02264_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_12054_ _06797_ VGND VGND VPWR VPWR _01546_ sky130_fd_sc_hd__clkbuf_1
X_16931_ clknet_leaf_8_clk _01257_ VGND VGND VPWR VPWR per_uart.uart0.txd_reg\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_11005_ net2290 _05719_ _06201_ VGND VGND VPWR VPWR _06205_ sky130_fd_sc_hd__mux2_1
X_16862_ _04150_ VGND VGND VPWR VPWR _02624_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_144_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15813_ CPU.registerFile\[12\]\[12\] _03118_ VGND VGND VPWR VPWR _03300_ sky130_fd_sc_hd__or2_1
X_16793_ _05289_ _04945_ _07132_ VGND VGND VPWR VPWR _04104_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15744_ CPU.registerFile\[21\]\[10\] CPU.registerFile\[23\]\[10\] _05441_ VGND VGND
+ VPWR VPWR _03233_ sky130_fd_sc_hd__mux2_1
X_12956_ _07305_ VGND VGND VPWR VPWR _07397_ sky130_fd_sc_hd__buf_4
XFILLER_0_158_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11907_ _06719_ VGND VGND VPWR VPWR _01616_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_47_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13988__270 clknet_1_1__leaf__08359_ VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__inv_2
X_15675_ _02771_ _03163_ _03164_ _03165_ _02782_ VGND VGND VPWR VPWR _03166_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_16_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_250 _03663_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12887_ CPU.registerFile\[21\]\[1\] _07289_ _07290_ CPU.registerFile\[17\]\[1\] _07300_
+ VGND VGND VPWR VPWR _07329_ sky130_fd_sc_hd__o221a_1
XANTENNA_261 _05066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_272 _05528_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17414_ net603 _01702_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[7\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_283 _05594_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11838_ net1707 _05685_ _06675_ VGND VGND VPWR VPWR _06683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_294 _07271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17345_ net534 _01633_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[9\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_60_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11769_ _06646_ VGND VGND VPWR VPWR _01681_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13508_ CPU.registerFile\[6\]\[18\] CPU.registerFile\[7\]\[18\] _07371_ VGND VGND
+ VPWR VPWR _07933_ sky130_fd_sc_hd__mux2_1
X_17276_ net465 _01564_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_155_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16227_ CPU.registerFile\[15\]\[24\] CPU.registerFile\[11\]\[24\] _02906_ VGND VGND
+ VPWR VPWR _03702_ sky130_fd_sc_hd__mux2_1
X_13439_ _07653_ _07864_ _07865_ VGND VGND VPWR VPWR _07866_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_24_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16158_ _03633_ _03634_ _02875_ VGND VGND VPWR VPWR _03635_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15109_ _07193_ net1432 _02726_ VGND VGND VPWR VPWR _02284_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16089_ CPU.registerFile\[7\]\[20\] _02898_ _02999_ _03567_ VGND VGND VPWR VPWR _03568_
+ sky130_fd_sc_hd__o211a_1
X_08980_ _04213_ VGND VGND VPWR VPWR _04698_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_58_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09601_ _04277_ _04406_ _04422_ VGND VGND VPWR VPWR _05296_ sky130_fd_sc_hd__nor3_1
X_09532_ _05229_ VGND VGND VPWR VPWR _05230_ sky130_fd_sc_hd__buf_4
XFILLER_0_149_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09463_ CPU.aluReg\[12\] _04808_ _05157_ _05163_ VGND VGND VPWR VPWR _05164_ sky130_fd_sc_hd__a211o_1
XFILLER_0_19_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09394_ CPU.Jimm\[15\] _04498_ _04503_ CPU.cycles\[15\] _05097_ VGND VGND VPWR VPWR
+ _05098_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_788 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_126_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14644__753 clknet_1_0__leaf__02680_ VGND VGND VPWR VPWR net785 sky130_fd_sc_hd__inv_2
X_16636__81 clknet_1_1__leaf__03988_ VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__inv_2
X_12810_ _07252_ VGND VGND VPWR VPWR _07253_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13790_ CPU.registerFile\[2\]\[27\] _07621_ VGND VGND VPWR VPWR _08206_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_2_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14945__1024 clknet_1_1__leaf__02710_ VGND VGND VPWR VPWR net1056 sky130_fd_sc_hd__inv_2
X_12741_ per_uart.d_in_uart\[0\] _07177_ _07203_ per_uart.uart0.txd_reg\[1\] VGND
+ VGND VPWR VPWR _07217_ sky130_fd_sc_hd__a22o_1
X_16651__95 clknet_1_0__leaf__03989_ VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__inv_2
XFILLER_0_38_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15460_ _02935_ _02947_ _02956_ _07703_ VGND VGND VPWR VPWR _02957_ sky130_fd_sc_hd__a31o_1
X_12672_ net1491 _07162_ VGND VGND VPWR VPWR _00029_ sky130_fd_sc_hd__xor2_1
XFILLER_0_155_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11623_ mapped_spi_ram.snd_bitcount\[5\] _06551_ VGND VGND VPWR VPWR _06553_ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15391_ _02791_ VGND VGND VPWR VPWR _02889_ sky130_fd_sc_hd__buf_4
X_14042__319 clknet_1_1__leaf__08364_ VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__inv_2
XFILLER_0_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_22_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_8
X_17130_ clknet_leaf_22_clk _00033_ VGND VGND VPWR VPWR CPU.cycles\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11554_ net1394 _06495_ _06505_ _06006_ VGND VGND VPWR VPWR _01754_ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17061_ net319 _01383_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_10505_ _05886_ _05911_ VGND VGND VPWR VPWR _05912_ sky130_fd_sc_hd__nor2_1
X_14273_ _04291_ net24 VGND VGND VPWR VPWR _08452_ sky130_fd_sc_hd__nand2_1
X_14690__795 clknet_1_0__leaf__02684_ VGND VGND VPWR VPWR net827 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_21_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11485_ _05541_ net2464 _06455_ VGND VGND VPWR VPWR _06460_ sky130_fd_sc_hd__mux2_1
X_16012_ CPU.registerFile\[30\]\[17\] _05050_ _02923_ _03493_ VGND VGND VPWR VPWR
+ _03494_ sky130_fd_sc_hd__o211a_1
X_13224_ _07647_ _07657_ _07395_ VGND VGND VPWR VPWR _07658_ sky130_fd_sc_hd__o21a_1
Xclkbuf_0__02750_ _02750_ VGND VGND VPWR VPWR clknet_0__02750_ sky130_fd_sc_hd__clkbuf_16
X_10436_ net1385 _05849_ _05854_ _05855_ VGND VGND VPWR VPWR _02225_ sky130_fd_sc_hd__o211a_1
XFILLER_0_21_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__02681_ _02681_ VGND VGND VPWR VPWR clknet_0__02681_ sky130_fd_sc_hd__clkbuf_16
X_13155_ CPU.registerFile\[31\]\[7\] _07482_ _07420_ CPU.registerFile\[27\]\[7\] _07483_
+ VGND VGND VPWR VPWR _07591_ sky130_fd_sc_hd__o221a_1
X_10367_ _05805_ VGND VGND VPWR VPWR _02245_ sky130_fd_sc_hd__clkbuf_1
X_12106_ _04762_ net2092 _06819_ VGND VGND VPWR VPWR _06825_ sky130_fd_sc_hd__mux2_1
X_10298_ _05768_ VGND VGND VPWR VPWR _02292_ sky130_fd_sc_hd__clkbuf_1
X_17963_ net1151 _02247_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[8\] sky130_fd_sc_hd__dfxtp_1
X_14727__828 clknet_1_1__leaf__02688_ VGND VGND VPWR VPWR net860 sky130_fd_sc_hd__inv_2
X_13086_ CPU.registerFile\[30\]\[5\] CPU.registerFile\[26\]\[5\] _07297_ VGND VGND
+ VPWR VPWR _07524_ sky130_fd_sc_hd__mux2_1
X_12037_ _06788_ VGND VGND VPWR VPWR _01554_ sky130_fd_sc_hd__clkbuf_1
X_16914_ net1974 _04182_ VGND VGND VPWR VPWR _04186_ sky130_fd_sc_hd__or2_1
X_17894_ net1083 _02178_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16845_ net1540 per_uart.rx_data\[1\] _04139_ VGND VGND VPWR VPWR _04141_ sky130_fd_sc_hd__mux2_1
X_16776_ _04050_ _04087_ _04088_ _04089_ VGND VGND VPWR VPWR _04090_ sky130_fd_sc_hd__a31o_1
XFILLER_0_87_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15727_ CPU.registerFile\[22\]\[9\] _08399_ VGND VGND VPWR VPWR _03217_ sky130_fd_sc_hd__and2_1
X_12939_ _07379_ VGND VGND VPWR VPWR _07380_ sky130_fd_sc_hd__buf_4
XFILLER_0_158_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15658_ CPU.registerFile\[20\]\[7\] CPU.registerFile\[21\]\[7\] _03066_ VGND VGND
+ VPWR VPWR _03150_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_157_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_157_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15589_ _02760_ VGND VGND VPWR VPWR _03082_ sky130_fd_sc_hd__buf_4
Xclkbuf_leaf_13_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17328_ net517 _01616_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[24\] sky130_fd_sc_hd__dfxtp_1
Xclkbuf_1_1__f__03966_ clknet_0__03966_ VGND VGND VPWR VPWR clknet_1_1__leaf__03966_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_44_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17259_ net449 _01547_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_256 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08963_ _04504_ _04483_ _04208_ VGND VGND VPWR VPWR _04682_ sky130_fd_sc_hd__nand3_2
XFILLER_0_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08894_ _04594_ _04599_ _04613_ VGND VGND VPWR VPWR _04614_ sky130_fd_sc_hd__nor3_4
X_14366__503 clknet_1_0__leaf__02652_ VGND VGND VPWR VPWR net535 sky130_fd_sc_hd__inv_2
XFILLER_0_79_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__02670_ clknet_0__02670_ VGND VGND VPWR VPWR clknet_1_0__leaf__02670_
+ sky130_fd_sc_hd__clkbuf_16
X_09515_ _04776_ _05212_ _04636_ VGND VGND VPWR VPWR _05213_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_88_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_104_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09446_ _05142_ _05147_ _04492_ VGND VGND VPWR VPWR _05148_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_148_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09377_ _04333_ _04701_ _05081_ _04678_ VGND VGND VPWR VPWR _05082_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_148_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11270_ _06345_ VGND VGND VPWR VPWR _01882_ sky130_fd_sc_hd__clkbuf_1
X_10221_ net1978 _05723_ _05713_ VGND VGND VPWR VPWR _05724_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_18_Left_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10152_ _04730_ VGND VGND VPWR VPWR _05677_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_7_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10083_ _05638_ VGND VGND VPWR VPWR _02377_ sky130_fd_sc_hd__clkbuf_1
X_13911_ _07394_ _08309_ _08323_ _08015_ VGND VGND VPWR VPWR _08324_ sky130_fd_sc_hd__a211o_1
XFILLER_0_89_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13842_ CPU.registerFile\[5\]\[28\] CPU.registerFile\[4\]\[28\] _04986_ VGND VGND
+ VPWR VPWR _08257_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13773_ CPU.registerFile\[28\]\[26\] CPU.registerFile\[24\]\[26\] _07476_ VGND VGND
+ VPWR VPWR _08190_ sky130_fd_sc_hd__mux2_1
X_10985_ _06194_ VGND VGND VPWR VPWR _02016_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_27_Left_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15512_ CPU.registerFile\[6\]\[4\] CPU.registerFile\[7\]\[4\] _02870_ VGND VGND VPWR
+ VPWR _03007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18300_ net34 _02580_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_12724_ _07204_ net1587 _07205_ VGND VGND VPWR VPWR _07206_ sky130_fd_sc_hd__mux2_1
X_16492_ _03955_ _03959_ _02810_ VGND VGND VPWR VPWR _03960_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18231_ net72 _02511_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_15443_ _02779_ VGND VGND VPWR VPWR _02940_ sky130_fd_sc_hd__clkbuf_8
X_12655_ CPU.cycles\[15\] _07152_ VGND VGND VPWR VPWR _07154_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_139_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18162_ clknet_leaf_29_clk _02442_ VGND VGND VPWR VPWR CPU.aluIn1\[28\] sky130_fd_sc_hd__dfxtp_2
X_11606_ net1376 _06501_ _06496_ CPU.mem_wdata\[5\] _06508_ VGND VGND VPWR VPWR _06542_
+ sky130_fd_sc_hd__a221o_1
X_15374_ _02821_ VGND VGND VPWR VPWR _02872_ sky130_fd_sc_hd__buf_4
XFILLER_0_136_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12586_ _07116_ VGND VGND VPWR VPWR _01266_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15149__1177 clknet_1_1__leaf__02745_ VGND VGND VPWR VPWR net1209 sky130_fd_sc_hd__inv_2
X_17113_ clknet_leaf_18_clk _00046_ VGND VGND VPWR VPWR CPU.cycles\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18093_ net156 _02373_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_11537_ mapped_spi_ram.state\[1\] VGND VGND VPWR VPWR _06493_ sky130_fd_sc_hd__buf_2
XFILLER_0_151_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__02702_ clknet_0__02702_ VGND VGND VPWR VPWR clknet_1_1__leaf__02702_
+ sky130_fd_sc_hd__clkbuf_16
X_17044_ net302 _01366_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[6\] sky130_fd_sc_hd__dfxtp_1
Xhold409 CPU.registerFile\[28\]\[29\] VGND VGND VPWR VPWR net1650 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11468_ _05524_ net2532 _06444_ VGND VGND VPWR VPWR _06451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Left_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13207_ _07311_ VGND VGND VPWR VPWR _07641_ sky130_fd_sc_hd__buf_4
X_10419_ _04192_ VGND VGND VPWR VPWR _05843_ sky130_fd_sc_hd__buf_4
X_11399_ _06414_ VGND VGND VPWR VPWR _01822_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_55_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14315__457 clknet_1_1__leaf__08464_ VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_55_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _07570_ _07573_ VGND VGND VPWR VPWR _07574_ sky130_fd_sc_hd__or2_1
Xclkbuf_0__02664_ _02664_ VGND VGND VPWR VPWR clknet_0__02664_ sky130_fd_sc_hd__clkbuf_16
X_13953__239 clknet_1_1__leaf__07226_ VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__inv_2
X_17946_ net1135 _02230_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[26\] sky130_fd_sc_hd__dfxtp_1
X_13069_ _07499_ _07501_ _07504_ _07506_ VGND VGND VPWR VPWR _07507_ sky130_fd_sc_hd__a22o_2
Xhold1109 CPU.registerFile\[20\]\[8\] VGND VGND VPWR VPWR net2350 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_119_Right_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17877_ net1066 _02161_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_bitcount\[2\] sky130_fd_sc_hd__dfxtp_1
X_16828_ per_uart.uart0.tx_bitcount\[3\] _04128_ per_uart.uart0.tx_bitcount\[0\] VGND
+ VGND VPWR VPWR _04129_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_136_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16759_ _04071_ _04075_ _04015_ VGND VGND VPWR VPWR _02596_ sky130_fd_sc_hd__a21oi_1
X_09300_ net1719 _05008_ _04983_ VGND VGND VPWR VPWR _05009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16630__76 clknet_1_0__leaf__03971_ VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__inv_2
XFILLER_0_152_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14361__499 clknet_1_0__leaf__08468_ VGND VGND VPWR VPWR net531 sky130_fd_sc_hd__inv_2
X_09231_ CPU.aluIn1\[22\] _04239_ _04210_ VGND VGND VPWR VPWR _04942_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09162_ CPU.PC\[2\] _04870_ VGND VGND VPWR VPWR _04874_ sky130_fd_sc_hd__or2_1
XFILLER_0_145_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_882 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09093_ _04800_ _04802_ _04804_ _04678_ VGND VGND VPWR VPWR _04805_ sky130_fd_sc_hd__o211a_1
XFILLER_0_43_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold910 CPU.registerFile\[19\]\[2\] VGND VGND VPWR VPWR net2151 sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 CPU.registerFile\[29\]\[5\] VGND VGND VPWR VPWR net2162 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold932 CPU.registerFile\[12\]\[5\] VGND VGND VPWR VPWR net2173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold943 CPU.registerFile\[3\]\[20\] VGND VGND VPWR VPWR net2184 sky130_fd_sc_hd__dlygate4sd3_1
X_14944__1023 clknet_1_0__leaf__02710_ VGND VGND VPWR VPWR net1055 sky130_fd_sc_hd__inv_2
Xhold954 CPU.registerFile\[17\]\[25\] VGND VGND VPWR VPWR net2195 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold965 CPU.registerFile\[25\]\[18\] VGND VGND VPWR VPWR net2206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold976 CPU.registerFile\[7\]\[3\] VGND VGND VPWR VPWR net2217 sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 CPU.registerFile\[29\]\[27\] VGND VGND VPWR VPWR net2228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 CPU.registerFile\[17\]\[9\] VGND VGND VPWR VPWR net2239 sky130_fd_sc_hd__dlygate4sd3_1
X_09995_ _05590_ VGND VGND VPWR VPWR _02449_ sky130_fd_sc_hd__clkbuf_1
X_14071__345 clknet_1_0__leaf__08367_ VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_4_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08946_ _04663_ _04664_ CPU.writeBack _04665_ VGND VGND VPWR VPWR _04666_ sky130_fd_sc_hd__or4bb_4
XTAP_TAPCELL_ROW_4_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08877_ _04578_ _04595_ VGND VGND VPWR VPWR _04597_ sky130_fd_sc_hd__or2_1
Xclkbuf_1_0__f__02722_ clknet_0__02722_ VGND VGND VPWR VPWR clknet_1_0__leaf__02722_
+ sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0__f__02653_ clknet_0__02653_ VGND VGND VPWR VPWR clknet_1_0__leaf__02653_
+ sky130_fd_sc_hd__clkbuf_16
X_10770_ _05509_ net2001 _06070_ VGND VGND VPWR VPWR _06080_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14756__854 clknet_1_0__leaf__02691_ VGND VGND VPWR VPWR net886 sky130_fd_sc_hd__inv_2
X_09429_ _05131_ VGND VGND VPWR VPWR _02564_ sky130_fd_sc_hd__clkbuf_1
X_12440_ _07039_ VGND VGND VPWR VPWR _01368_ sky130_fd_sc_hd__clkbuf_1
X_16516__184 clknet_1_0__leaf__03963_ VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__inv_2
XFILLER_0_34_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12371_ _05253_ net1901 _06999_ VGND VGND VPWR VPWR _07003_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14110_ _08383_ VGND VGND VPWR VPWR _01464_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_134_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11322_ _06373_ VGND VGND VPWR VPWR _01858_ sky130_fd_sc_hd__clkbuf_1
X_15090_ net1423 _07182_ net1464 VGND VGND VPWR VPWR _02732_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_105_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11253_ CPU.registerFile\[9\]\[20\] _05694_ _06335_ VGND VGND VPWR VPWR _06337_ sky130_fd_sc_hd__mux2_1
X_10204_ _05187_ VGND VGND VPWR VPWR _05712_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11184_ _06300_ VGND VGND VPWR VPWR _01923_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17800_ net989 _02084_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_10135_ _05665_ VGND VGND VPWR VPWR _02352_ sky130_fd_sc_hd__clkbuf_1
X_15992_ CPU.registerFile\[16\]\[17\] CPU.registerFile\[18\]\[17\] _03032_ VGND VGND
+ VPWR VPWR _03474_ sky130_fd_sc_hd__mux2_1
X_17731_ net920 _02015_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_10066_ _05628_ VGND VGND VPWR VPWR _02384_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_50_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03969_ clknet_0__03969_ VGND VGND VPWR VPWR clknet_1_0__leaf__03969_
+ sky130_fd_sc_hd__clkbuf_16
X_17662_ net851 _01950_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13825_ CPU.registerFile\[15\]\[28\] _07772_ _07773_ CPU.registerFile\[11\]\[28\]
+ _08239_ VGND VGND VPWR VPWR _08240_ sky130_fd_sc_hd__o221a_1
X_16613_ net1552 net2069 _03979_ VGND VGND VPWR VPWR _03982_ sky130_fd_sc_hd__mux2_1
X_17593_ net782 _01881_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[11\] sky130_fd_sc_hd__dfxtp_1
X_14839__929 clknet_1_0__leaf__02699_ VGND VGND VPWR VPWR net961 sky130_fd_sc_hd__inv_2
XFILLER_0_58_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16544_ clknet_1_0__leaf__07219_ VGND VGND VPWR VPWR _03966_ sky130_fd_sc_hd__buf_1
XFILLER_0_15_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13756_ _07380_ _08165_ _08173_ _07703_ VGND VGND VPWR VPWR _08174_ sky130_fd_sc_hd__a31o_1
X_10968_ _06185_ VGND VGND VPWR VPWR _02024_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__08358_ clknet_0__08358_ VGND VGND VPWR VPWR clknet_1_0__leaf__08358_
+ sky130_fd_sc_hd__clkbuf_16
X_12707_ net1457 _07188_ VGND VGND VPWR VPWR _07189_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16475_ CPU.registerFile\[8\]\[31\] CPU.registerFile\[12\]\[31\] _03254_ VGND VGND
+ VPWR VPWR _03943_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13687_ CPU.registerFile\[13\]\[23\] _07403_ _07404_ CPU.registerFile\[9\]\[23\]
+ _07250_ VGND VGND VPWR VPWR _08107_ sky130_fd_sc_hd__o221a_1
X_10899_ net1599 _05681_ _06143_ VGND VGND VPWR VPWR _06149_ sky130_fd_sc_hd__mux2_1
X_18214_ net55 _02494_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_15426_ _02769_ VGND VGND VPWR VPWR _02923_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12638_ CPU.cycles\[7\] CPU.cycles\[8\] _07142_ VGND VGND VPWR VPWR _07144_ sky130_fd_sc_hd__and3_1
X_16928__8 clknet_1_1__leaf__07220_ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__inv_2
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18145_ clknet_leaf_19_clk _02425_ VGND VGND VPWR VPWR CPU.aluIn1\[11\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_124_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15357_ _02854_ VGND VGND VPWR VPWR _02855_ sky130_fd_sc_hd__clkbuf_8
X_12569_ CPU.registerFile\[4\]\[11\] _05187_ _07107_ VGND VGND VPWR VPWR _07108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_44_Left_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18076_ net139 _02356_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_15288_ _02760_ VGND VGND VPWR VPWR _02787_ sky130_fd_sc_hd__clkbuf_8
Xhold206 CPU.cycles\[24\] VGND VGND VPWR VPWR net1447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold217 mapped_spi_flash.rcv_data\[18\] VGND VGND VPWR VPWR net1458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 _02193_ VGND VGND VPWR VPWR net1469 sky130_fd_sc_hd__dlygate4sd3_1
X_17027_ net285 _01349_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold239 CPU.rs2\[24\] VGND VGND VPWR VPWR net1480 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0__02716_ _02716_ VGND VGND VPWR VPWR clknet_0__02716_ sky130_fd_sc_hd__clkbuf_16
X_15222__132 clknet_1_1__leaf__02753_ VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__inv_2
XFILLER_0_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08800_ _04518_ _04519_ VGND VGND VPWR VPWR _04520_ sky130_fd_sc_hd__and2_4
X_09780_ _05460_ VGND VGND VPWR VPWR _02534_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08731_ _04450_ VGND VGND VPWR VPWR _04451_ sky130_fd_sc_hd__inv_2
X_17929_ net1118 _02213_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[9\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_53_Left_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08662_ _04381_ _04237_ VGND VGND VPWR VPWR _04382_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_68_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08593_ CPU.aluIn1\[7\] _04272_ VGND VGND VPWR VPWR _04313_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14478__604 clknet_1_1__leaf__02663_ VGND VGND VPWR VPWR net636 sky130_fd_sc_hd__inv_2
XFILLER_0_9_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09214_ CPU.PC\[17\] _04925_ VGND VGND VPWR VPWR _04926_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_62_Left_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_901 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09145_ CPU.PC\[10\] CPU.Bimm\[10\] _04820_ VGND VGND VPWR VPWR _04857_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09076_ _04238_ _04347_ _04348_ VGND VGND VPWR VPWR _04789_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_116_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold740 CPU.registerFile\[31\]\[3\] VGND VGND VPWR VPWR net1981 sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 CPU.registerFile\[23\]\[27\] VGND VGND VPWR VPWR net1992 sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 CPU.registerFile\[1\]\[10\] VGND VGND VPWR VPWR net2003 sky130_fd_sc_hd__dlygate4sd3_1
Xhold773 CPU.registerFile\[20\]\[12\] VGND VGND VPWR VPWR net2014 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_899 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold784 CPU.registerFile\[15\]\[1\] VGND VGND VPWR VPWR net2025 sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 CPU.registerFile\[13\]\[10\] VGND VGND VPWR VPWR net2036 sky130_fd_sc_hd__dlygate4sd3_1
X_09978_ _05532_ net1880 _05581_ VGND VGND VPWR VPWR _05582_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_71_Left_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08929_ _04647_ _04648_ _04621_ VGND VGND VPWR VPWR _04649_ sky130_fd_sc_hd__mux2_4
X_15148__1176 clknet_1_1__leaf__02745_ VGND VGND VPWR VPWR net1208 sky130_fd_sc_hd__inv_2
X_11940_ net2447 _05719_ _06733_ VGND VGND VPWR VPWR _06737_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11871_ _06700_ VGND VGND VPWR VPWR _01633_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__02705_ clknet_0__02705_ VGND VGND VPWR VPWR clknet_1_0__leaf__02705_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_98_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13610_ _08028_ _08031_ _07405_ VGND VGND VPWR VPWR _08032_ sky130_fd_sc_hd__mux2_1
X_10822_ net1639 _05673_ _06106_ VGND VGND VPWR VPWR _06108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14344__483 clknet_1_0__leaf__08467_ VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__inv_2
X_13541_ CPU.registerFile\[2\]\[19\] _07388_ VGND VGND VPWR VPWR _07965_ sky130_fd_sc_hd__or2_1
X_10753_ _06071_ VGND VGND VPWR VPWR _02125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16260_ _02812_ _03731_ _03733_ _02767_ VGND VGND VPWR VPWR _03734_ sky130_fd_sc_hd__a211o_1
X_13982__265 clknet_1_0__leaf__08358_ VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__inv_2
X_13472_ CPU.registerFile\[31\]\[17\] _07382_ _07383_ CPU.registerFile\[27\]\[17\]
+ _07254_ VGND VGND VPWR VPWR _07898_ sky130_fd_sc_hd__o221a_1
X_10684_ _05487_ CPU.registerFile\[28\]\[31\] _06034_ VGND VGND VPWR VPWR _06035_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12423_ _07030_ VGND VGND VPWR VPWR _01376_ sky130_fd_sc_hd__clkbuf_1
X_16191_ CPU.registerFile\[1\]\[23\] _02822_ _03666_ _02887_ VGND VGND VPWR VPWR _03667_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12354_ _05090_ net1863 _06988_ VGND VGND VPWR VPWR _06994_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11305_ _06364_ VGND VGND VPWR VPWR _01866_ sky130_fd_sc_hd__clkbuf_1
X_12285_ CPU.aluReg\[9\] CPU.aluReg\[7\] _06939_ VGND VGND VPWR VPWR _06949_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11236_ net2453 _05677_ _06324_ VGND VGND VPWR VPWR _06328_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11167_ _06291_ VGND VGND VPWR VPWR _01931_ sky130_fd_sc_hd__clkbuf_1
X_10118_ net2306 _05209_ _05655_ VGND VGND VPWR VPWR _05657_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_147_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11098_ net2047 _05675_ _06252_ VGND VGND VPWR VPWR _06255_ sky130_fd_sc_hd__mux2_1
X_15975_ CPU.registerFile\[22\]\[16\] CPU.registerFile\[23\]\[16\] _02828_ VGND VGND
+ VPWR VPWR _03458_ sky130_fd_sc_hd__mux2_1
X_17714_ net903 _01998_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10049_ net2364 _05209_ _05618_ VGND VGND VPWR VPWR _05620_ sky130_fd_sc_hd__mux2_1
X_14427__558 clknet_1_1__leaf__02658_ VGND VGND VPWR VPWR net590 sky130_fd_sc_hd__inv_2
X_17645_ net834 _01933_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13808_ CPU.registerFile\[9\]\[27\] _07618_ _08223_ _07417_ _07554_ VGND VGND VPWR
+ VPWR _08224_ sky130_fd_sc_hd__o221a_1
X_17576_ net765 _01864_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14943__1022 clknet_1_1__leaf__02710_ VGND VGND VPWR VPWR net1054 sky130_fd_sc_hd__inv_2
XFILLER_0_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13739_ _04814_ _08152_ _08156_ _07271_ VGND VGND VPWR VPWR _08157_ sky130_fd_sc_hd__a211o_1
XFILLER_0_128_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16458_ _08411_ _03919_ _03926_ _07308_ VGND VGND VPWR VPWR _03927_ sky130_fd_sc_hd__a31o_1
XFILLER_0_144_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15409_ _02772_ VGND VGND VPWR VPWR _02906_ sky130_fd_sc_hd__buf_4
XFILLER_0_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16389_ _03856_ _03859_ _02809_ VGND VGND VPWR VPWR _03860_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18128_ net191 _02408_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[26\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_124_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18059_ net1232 _02339_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09901_ _05535_ net2168 _05533_ VGND VGND VPWR VPWR _05536_ sky130_fd_sc_hd__mux2_1
XFILLER_0_158_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14785__880 clknet_1_0__leaf__02694_ VGND VGND VPWR VPWR net912 sky130_fd_sc_hd__inv_2
X_09832_ _04660_ _04661_ VGND VGND VPWR VPWR _05488_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_111_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09763_ _04666_ _05450_ VGND VGND VPWR VPWR _05451_ sky130_fd_sc_hd__nor2_2
X_08714_ _04400_ _04430_ _04401_ _04431_ _04433_ VGND VGND VPWR VPWR _04434_ sky130_fd_sc_hd__o311a_4
X_09694_ mapped_spi_ram.rcv_data\[26\] net17 net1290 per_uart.rx_data\[2\] VGND VGND
+ VPWR VPWR _05385_ sky130_fd_sc_hd__a22o_1
Xrebuffer10 net1252 VGND VGND VPWR VPWR net1251 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer21 net1263 VGND VGND VPWR VPWR net1262 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer32 net1272 VGND VGND VPWR VPWR net1273 sky130_fd_sc_hd__dlygate4sd1_1
X_08645_ _04226_ _04364_ VGND VGND VPWR VPWR _04365_ sky130_fd_sc_hd__and2b_1
Xrebuffer43 net1286 VGND VGND VPWR VPWR net1284 sky130_fd_sc_hd__buf_2
XFILLER_0_49_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08576_ CPU.Iimm\[1\] VGND VGND VPWR VPWR _04296_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_138_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_864 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_845 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_558 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09128_ CPU.PC\[17\] _04838_ VGND VGND VPWR VPWR _04840_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_98_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14868__955 clknet_1_1__leaf__02702_ VGND VGND VPWR VPWR net987 sky130_fd_sc_hd__inv_2
X_09059_ _04491_ VGND VGND VPWR VPWR _04773_ sky130_fd_sc_hd__clkbuf_4
X_12070_ _05188_ net2052 _06805_ VGND VGND VPWR VPWR _06806_ sky130_fd_sc_hd__mux2_1
Xhold570 CPU.registerFile\[29\]\[22\] VGND VGND VPWR VPWR net1811 sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 CPU.registerFile\[2\]\[21\] VGND VGND VPWR VPWR net1822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 CPU.registerFile\[7\]\[11\] VGND VGND VPWR VPWR net1833 sky130_fd_sc_hd__dlygate4sd3_1
X_11021_ net1589 _05735_ _06178_ VGND VGND VPWR VPWR _06213_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15760_ CPU.registerFile\[9\]\[10\] _08404_ _05071_ VGND VGND VPWR VPWR _03249_ sky130_fd_sc_hd__o21a_1
X_12972_ CPU.registerFile\[14\]\[2\] CPU.registerFile\[10\]\[2\] _07399_ VGND VGND
+ VPWR VPWR _07413_ sky130_fd_sc_hd__mux2_1
Xhold1270 CPU.registerFile\[15\]\[9\] VGND VGND VPWR VPWR net2511 sky130_fd_sc_hd__dlygate4sd3_1
X_11923_ CPU.registerFile\[11\]\[16\] _05702_ _06722_ VGND VGND VPWR VPWR _06728_
+ sky130_fd_sc_hd__mux2_1
Xhold1281 CPU.aluReg\[2\] VGND VGND VPWR VPWR net2522 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15691_ _02812_ _03178_ _03181_ _02948_ VGND VGND VPWR VPWR _03182_ sky130_fd_sc_hd__o211a_1
Xhold1292 mapped_spi_flash.rcv_data\[14\] VGND VGND VPWR VPWR net2533 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_410 _04659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17430_ net619 _01718_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[23\] sky130_fd_sc_hd__dfxtp_1
X_11854_ _06691_ VGND VGND VPWR VPWR _01641_ sky130_fd_sc_hd__clkbuf_1
X_10805_ _06098_ VGND VGND VPWR VPWR _02100_ sky130_fd_sc_hd__clkbuf_1
X_17361_ net550 _01649_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_14573_ clknet_1_0__leaf__02664_ VGND VGND VPWR VPWR _02673_ sky130_fd_sc_hd__buf_1
X_11785_ net1244 net1914 _06650_ VGND VGND VPWR VPWR _06655_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13524_ CPU.registerFile\[28\]\[18\] CPU.registerFile\[24\]\[18\] _07492_ VGND VGND
+ VPWR VPWR _07949_ sky130_fd_sc_hd__mux2_1
X_16312_ _02856_ _03782_ _03784_ _02794_ VGND VGND VPWR VPWR _03785_ sky130_fd_sc_hd__o211a_1
X_17292_ net481 _01580_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_10736_ _05543_ net2200 _06056_ VGND VGND VPWR VPWR _06062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_137_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16243_ CPU.registerFile\[2\]\[24\] _03143_ _02822_ CPU.registerFile\[3\]\[24\] _03144_
+ VGND VGND VPWR VPWR _03718_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_11_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13455_ CPU.registerFile\[30\]\[16\] CPU.registerFile\[26\]\[16\] _04937_ VGND VGND
+ VPWR VPWR _07882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10667_ net1522 _06018_ _06022_ _06023_ VGND VGND VPWR VPWR _02163_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12406_ _07021_ VGND VGND VPWR VPWR _01384_ sky130_fd_sc_hd__clkbuf_1
X_16174_ CPU.registerFile\[20\]\[22\] CPU.registerFile\[21\]\[22\] _08395_ VGND VGND
+ VPWR VPWR _03651_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13386_ _07650_ _07813_ _07814_ VGND VGND VPWR VPWR _07815_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_112_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10598_ _05969_ VGND VGND VPWR VPWR _05981_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_152_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12337_ _04798_ net1728 _06977_ VGND VGND VPWR VPWR _06985_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_149_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12268_ CPU.aluReg\[13\] CPU.aluReg\[11\] _06906_ VGND VGND VPWR VPWR _06936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11219_ _06318_ VGND VGND VPWR VPWR _01906_ sky130_fd_sc_hd__clkbuf_1
X_12199_ CPU.aluReg\[29\] CPU.aluReg\[27\] _06871_ VGND VGND VPWR VPWR _06883_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15958_ CPU.registerFile\[28\]\[16\] _03064_ VGND VGND VPWR VPWR _03441_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_606 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15889_ _03369_ _03373_ _08410_ VGND VGND VPWR VPWR _03374_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_65_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17628_ net817 _01916_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17559_ net748 _01847_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_720 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15147__1175 clknet_1_1__leaf__02745_ VGND VGND VPWR VPWR net1207 sky130_fd_sc_hd__inv_2
XFILLER_0_6_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09815_ net2282 _05273_ _05474_ VGND VGND VPWR VPWR _05479_ sky130_fd_sc_hd__mux2_1
X_09746_ _05432_ _04481_ VGND VGND VPWR VPWR _05435_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09677_ _05368_ _04417_ VGND VGND VPWR VPWR _05369_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_38_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08628_ CPU.aluIn1\[23\] _04237_ VGND VGND VPWR VPWR _04348_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_124_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08559_ CPU.mem_wdata\[5\] CPU.Bimm\[5\] _04203_ VGND VGND VPWR VPWR _04279_ sky130_fd_sc_hd__mux2_2
XFILLER_0_37_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_823 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11570_ _06512_ _05895_ VGND VGND VPWR VPWR _06518_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10521_ net1384 _05892_ _05925_ _05885_ VGND VGND VPWR VPWR _02210_ sky130_fd_sc_hd__o211a_1
X_13240_ net2448 _07358_ _07658_ _07673_ _05844_ VGND VGND VPWR VPWR _01304_ sky130_fd_sc_hd__o221a_1
X_10452_ net1365 _05849_ _05866_ _05855_ VGND VGND VPWR VPWR _02220_ sky130_fd_sc_hd__o211a_1
X_14456__584 clknet_1_1__leaf__02661_ VGND VGND VPWR VPWR net616 sky130_fd_sc_hd__inv_2
X_13171_ _07245_ _07605_ VGND VGND VPWR VPWR _07606_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10383_ _04589_ VGND VGND VPWR VPWR _05815_ sky130_fd_sc_hd__buf_4
X_14194__372 clknet_1_1__leaf__08429_ VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__inv_2
X_12122_ _06833_ VGND VGND VPWR VPWR _01514_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14942__1021 clknet_1_0__leaf__02710_ VGND VGND VPWR VPWR net1053 sky130_fd_sc_hd__inv_2
X_12053_ _05027_ net1875 _06794_ VGND VGND VPWR VPWR _06797_ sky130_fd_sc_hd__mux2_1
X_16930_ clknet_leaf_8_clk _01256_ VGND VGND VPWR VPWR per_uart.uart0.txd_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_11004_ _06204_ VGND VGND VPWR VPWR _02007_ sky130_fd_sc_hd__clkbuf_1
X_16861_ _04138_ _04149_ _04193_ VGND VGND VPWR VPWR _04150_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_144_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15812_ CPU.registerFile\[14\]\[12\] CPU.registerFile\[10\]\[12\] _03082_ VGND VGND
+ VPWR VPWR _03299_ sky130_fd_sc_hd__mux2_1
X_16792_ _04052_ _04954_ _08453_ VGND VGND VPWR VPWR _04103_ sky130_fd_sc_hd__or3b_1
X_15743_ _03226_ _03231_ _08401_ VGND VGND VPWR VPWR _03232_ sky130_fd_sc_hd__mux2_1
X_12955_ _07381_ _07393_ _07395_ VGND VGND VPWR VPWR _07396_ sky130_fd_sc_hd__o21a_1
X_14621__732 clknet_1_0__leaf__02678_ VGND VGND VPWR VPWR net764 sky130_fd_sc_hd__inv_2
X_11906_ net1991 _05685_ _06711_ VGND VGND VPWR VPWR _06719_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15674_ CPU.registerFile\[9\]\[8\] _02778_ _03125_ VGND VGND VPWR VPWR _03165_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_16_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_240 _03004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12886_ CPU.registerFile\[23\]\[1\] _07325_ _07326_ CPU.registerFile\[19\]\[1\] _07327_
+ VGND VGND VPWR VPWR _07328_ sky130_fd_sc_hd__o221a_1
XFILLER_0_87_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_251 _05026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_262 _05071_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17413_ net602 net1331 VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_273 _05530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11837_ _06682_ VGND VGND VPWR VPWR _01649_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_284 _05594_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_295 _07271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17344_ net533 _01632_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_60_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ _04780_ net1792 _06639_ VGND VGND VPWR VPWR _06646_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_60_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14539__659 clknet_1_0__leaf__02669_ VGND VGND VPWR VPWR net691 sky130_fd_sc_hd__inv_2
XFILLER_0_126_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13507_ CPU.registerFile\[1\]\[18\] _07576_ _07931_ _07639_ VGND VGND VPWR VPWR _07932_
+ sky130_fd_sc_hd__a22o_1
X_10719_ _05526_ net1670 _06045_ VGND VGND VPWR VPWR _06053_ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17275_ net464 _01563_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_11699_ _06574_ VGND VGND VPWR VPWR _06603_ sky130_fd_sc_hd__buf_2
X_16226_ _02786_ _03698_ _03700_ _03019_ VGND VGND VPWR VPWR _03701_ sky130_fd_sc_hd__a211o_1
X_13438_ CPU.registerFile\[23\]\[16\] _07382_ _07383_ CPU.registerFile\[19\]\[16\]
+ _07288_ VGND VGND VPWR VPWR _07865_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_155_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer1 _04335_ VGND VGND VPWR VPWR net1242 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_23_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16157_ CPU.registerFile\[8\]\[22\] CPU.registerFile\[12\]\[22\] _08403_ VGND VGND
+ VPWR VPWR _03634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13369_ _07305_ _07788_ _07791_ _07232_ _07798_ VGND VGND VPWR VPWR _07799_ sky130_fd_sc_hd__o311a_2
X_15108_ per_uart.uart0.enable16_counter\[13\] _07191_ net1431 VGND VGND VPWR VPWR
+ _02741_ sky130_fd_sc_hd__o21ai_1
X_16088_ CPU.registerFile\[6\]\[20\] _02819_ VGND VGND VPWR VPWR _03567_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_58_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15039_ _02719_ VGND VGND VPWR VPWR _02236_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09600_ CPU.cycles\[6\] _04989_ _05290_ _05292_ _05294_ VGND VGND VPWR VPWR _05295_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14284__429 clknet_1_0__leaf__08435_ VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__inv_2
X_09531_ _05214_ _05223_ _05228_ VGND VGND VPWR VPWR _05229_ sky130_fd_sc_hd__or3b_4
X_15063__1129 clknet_1_1__leaf__02722_ VGND VGND VPWR VPWR net1161 sky130_fd_sc_hd__inv_2
XFILLER_0_79_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire23 _04191_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
X_14897__981 clknet_1_0__leaf__02705_ VGND VGND VPWR VPWR net1013 sky130_fd_sc_hd__inv_2
X_09462_ _04432_ _04488_ _05162_ _04677_ VGND VGND VPWR VPWR _05163_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09393_ _04817_ _05095_ _05096_ _04916_ VGND VGND VPWR VPWR _05097_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_47_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14750__849 clknet_1_1__leaf__02690_ VGND VGND VPWR VPWR net881 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_95_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16510__179 clknet_1_0__leaf__03962_ VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__inv_2
XFILLER_0_15_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_126_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09729_ _04672_ _05418_ VGND VGND VPWR VPWR _05419_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_2_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12740_ _07216_ VGND VGND VPWR VPWR _01261_ sky130_fd_sc_hd__clkbuf_1
X_12671_ _07162_ _07163_ VGND VGND VPWR VPWR _00028_ sky130_fd_sc_hd__nor2_1
X_11622_ mapped_spi_ram.snd_bitcount\[5\] _06551_ VGND VGND VPWR VPWR _06552_ sky130_fd_sc_hd__or2_1
X_15390_ CPU.registerFile\[31\]\[1\] _02887_ VGND VGND VPWR VPWR _02888_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11553_ net1389 _06499_ _06489_ _06504_ VGND VGND VPWR VPWR _06505_ sky130_fd_sc_hd__a211o_1
XFILLER_0_53_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17060_ net318 _01382_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_10504_ CPU.PC\[8\] _05867_ _05909_ _05910_ VGND VGND VPWR VPWR _05911_ sky130_fd_sc_hd__o2bb2a_4
X_14272_ _04701_ _08450_ _05435_ VGND VGND VPWR VPWR _08451_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11484_ _06459_ VGND VGND VPWR VPWR _01782_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_21_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16011_ CPU.registerFile\[26\]\[17\] _02861_ VGND VGND VPWR VPWR _03493_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13223_ _07652_ _07656_ _07584_ VGND VGND VPWR VPWR _07657_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_111_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10435_ _05843_ VGND VGND VPWR VPWR _05855_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0__02680_ _02680_ VGND VGND VPWR VPWR clknet_0__02680_ sky130_fd_sc_hd__clkbuf_16
X_13154_ CPU.registerFile\[30\]\[7\] CPU.registerFile\[26\]\[7\] _07480_ VGND VGND
+ VPWR VPWR _07590_ sky130_fd_sc_hd__mux2_1
X_10366_ _05543_ net2395 _05799_ VGND VGND VPWR VPWR _05805_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12105_ _06824_ VGND VGND VPWR VPWR _01522_ sky130_fd_sc_hd__clkbuf_1
X_17962_ net1150 _02246_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_13085_ _07519_ _07520_ _07522_ VGND VGND VPWR VPWR _07523_ sky130_fd_sc_hd__o21a_1
X_10297_ _05543_ net2202 _05762_ VGND VGND VPWR VPWR _05768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12036_ _04748_ net2285 _06783_ VGND VGND VPWR VPWR _06788_ sky130_fd_sc_hd__mux2_1
X_16913_ CPU.mem_wdata\[2\] _04180_ _04185_ _04176_ VGND VGND VPWR VPWR _02640_ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17893_ net1082 _02177_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[11\] sky130_fd_sc_hd__dfxtp_1
X_16844_ net1509 VGND VGND VPWR VPWR _02616_ sky130_fd_sc_hd__clkbuf_1
X_16775_ _04914_ _05015_ _03990_ VGND VGND VPWR VPWR _04089_ sky130_fd_sc_hd__a21o_1
X_15146__1174 clknet_1_0__leaf__02745_ VGND VGND VPWR VPWR net1206 sky130_fd_sc_hd__inv_2
X_13987_ clknet_1_0__leaf__07223_ VGND VGND VPWR VPWR _08359_ sky130_fd_sc_hd__buf_1
X_15726_ CPU.registerFile\[21\]\[9\] CPU.registerFile\[23\]\[9\] _02769_ VGND VGND
+ VPWR VPWR _03216_ sky130_fd_sc_hd__mux2_1
X_12938_ _07253_ VGND VGND VPWR VPWR _07379_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15657_ _03142_ _03145_ _03148_ _02945_ VGND VGND VPWR VPWR _03149_ sky130_fd_sc_hd__o22a_2
X_12869_ _05337_ VGND VGND VPWR VPWR _07311_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_157_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_157_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15588_ _07228_ VGND VGND VPWR VPWR _03081_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17327_ net516 _01615_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_1__f__03965_ clknet_0__03965_ VGND VGND VPWR VPWR clknet_1_1__leaf__03965_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_70_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17258_ net448 _01546_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_12_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16209_ CPU.registerFile\[9\]\[23\] CPU.registerFile\[13\]\[23\] _02851_ VGND VGND
+ VPWR VPWR _03685_ sky130_fd_sc_hd__mux2_1
X_17189_ clknet_leaf_25_clk _01477_ VGND VGND VPWR VPWR CPU.Jimm\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08962_ _04218_ VGND VGND VPWR VPWR _04681_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_90_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08893_ _04601_ _04604_ _04612_ VGND VGND VPWR VPWR _04613_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15191__104 clknet_1_1__leaf__02750_ VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__inv_2
XFILLER_0_78_200 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09514_ mapped_spi_ram.rcv_data\[17\] _04645_ _05211_ VGND VGND VPWR VPWR _05212_
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_88_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09445_ _04435_ _04806_ _05146_ _04679_ VGND VGND VPWR VPWR _05147_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_94_726 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_148_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_828 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14941__1020 clknet_1_0__leaf__02710_ VGND VGND VPWR VPWR net1052 sky130_fd_sc_hd__inv_2
XFILLER_0_148_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09376_ _05078_ _05080_ _04373_ VGND VGND VPWR VPWR _05081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10220_ _05305_ VGND VGND VPWR VPWR _05723_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10151_ _05676_ VGND VGND VPWR VPWR _02347_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10082_ net2317 _04748_ _05633_ VGND VGND VPWR VPWR _05638_ sky130_fd_sc_hd__mux2_1
X_14568__685 clknet_1_0__leaf__02672_ VGND VGND VPWR VPWR net717 sky130_fd_sc_hd__inv_2
X_13910_ _07334_ _08312_ _08315_ _08322_ _07766_ VGND VGND VPWR VPWR _08323_ sky130_fd_sc_hd__o311a_1
X_13841_ _08252_ _08255_ _07514_ VGND VGND VPWR VPWR _08256_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_69_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13772_ _08181_ _08188_ _07230_ VGND VGND VPWR VPWR _08189_ sky130_fd_sc_hd__o21a_1
X_10984_ net1765 _05698_ _06190_ VGND VGND VPWR VPWR _06194_ sky130_fd_sc_hd__mux2_1
X_15511_ CPU.registerFile\[1\]\[4\] _02867_ _03005_ _08405_ VGND VGND VPWR VPWR _03006_
+ sky130_fd_sc_hd__a22o_1
X_12723_ _07177_ _07203_ _04192_ VGND VGND VPWR VPWR _07205_ sky130_fd_sc_hd__o21ai_4
X_16491_ _02914_ _03956_ _03958_ _02864_ VGND VGND VPWR VPWR _03959_ sky130_fd_sc_hd__a211o_1
XFILLER_0_84_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18230_ net71 _02510_ VGND VGND VPWR VPWR CPU.registerFile\[19\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_15442_ _02813_ VGND VGND VPWR VPWR _02939_ sky130_fd_sc_hd__clkbuf_4
X_12654_ _07152_ net1488 VGND VGND VPWR VPWR _00020_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_139_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11605_ net1392 _06524_ _06541_ _06539_ VGND VGND VPWR VPWR _01739_ sky130_fd_sc_hd__o211a_1
X_18161_ clknet_leaf_29_clk _02441_ VGND VGND VPWR VPWR CPU.aluIn1\[27\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_81_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12585_ CPU.registerFile\[4\]\[3\] _05380_ _07107_ VGND VGND VPWR VPWR _07116_ sky130_fd_sc_hd__mux2_1
X_15373_ CPU.registerFile\[6\]\[1\] CPU.registerFile\[7\]\[1\] _02870_ VGND VGND VPWR
+ VPWR _02871_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14733__833 clknet_1_1__leaf__02689_ VGND VGND VPWR VPWR net865 sky130_fd_sc_hd__inv_2
X_17112_ clknet_leaf_23_clk _00045_ VGND VGND VPWR VPWR CPU.cycles\[8\] sky130_fd_sc_hd__dfxtp_1
X_11536_ _05816_ net1319 _06489_ _06492_ net1326 VGND VGND VPWR VPWR _01759_ sky130_fd_sc_hd__a32o_1
X_18092_ net155 _02372_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__02701_ clknet_0__02701_ VGND VGND VPWR VPWR clknet_1_1__leaf__02701_
+ sky130_fd_sc_hd__clkbuf_16
X_17043_ net301 _01365_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_11467_ _06450_ VGND VGND VPWR VPWR _01790_ sky130_fd_sc_hd__clkbuf_1
X_15062__1128 clknet_1_0__leaf__02722_ VGND VGND VPWR VPWR net1160 sky130_fd_sc_hd__inv_2
XFILLER_0_151_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13206_ CPU.registerFile\[1\]\[9\] _07576_ _07637_ _07639_ VGND VGND VPWR VPWR _07640_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10418_ mapped_spi_flash.state\[2\] _05817_ _05823_ VGND VGND VPWR VPWR _05842_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11398_ _05522_ net2305 _06408_ VGND VGND VPWR VPWR _06414_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_0__02663_ _02663_ VGND VGND VPWR VPWR clknet_0__02663_ sky130_fd_sc_hd__clkbuf_16
X_13137_ CPU.registerFile\[23\]\[7\] _07502_ _07503_ CPU.registerFile\[19\]\[7\] _07572_
+ VGND VGND VPWR VPWR _07573_ sky130_fd_sc_hd__o221a_1
X_10349_ _05526_ net2028 _05788_ VGND VGND VPWR VPWR _05796_ sky130_fd_sc_hd__mux2_1
X_17945_ net1134 _02229_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[25\] sky130_fd_sc_hd__dfxtp_1
X_13068_ _07330_ _07505_ VGND VGND VPWR VPWR _07506_ sky130_fd_sc_hd__or2_1
X_12019_ _06778_ VGND VGND VPWR VPWR _01563_ sky130_fd_sc_hd__clkbuf_1
X_17876_ net1065 _02160_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_bitcount\[1\] sky130_fd_sc_hd__dfxtp_1
X_16827_ per_uart.uart0.tx_bitcount\[2\] VGND VGND VPWR VPWR _04128_ sky130_fd_sc_hd__inv_2
X_16758_ _04050_ _04072_ _04073_ _04074_ VGND VGND VPWR VPWR _04075_ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15709_ _03195_ _03196_ _03198_ _02965_ VGND VGND VPWR VPWR _03199_ sky130_fd_sc_hd__a211o_1
XFILLER_0_75_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16689_ _07123_ _05291_ VGND VGND VPWR VPWR _04016_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09230_ CPU.Iimm\[2\] _04812_ _04503_ CPU.cycles\[22\] VGND VGND VPWR VPWR _04941_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14025__304 clknet_1_1__leaf__08362_ VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__inv_2
XFILLER_0_152_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09161_ CPU.PC\[1\] _04872_ VGND VGND VPWR VPWR _04873_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18359_ clknet_leaf_4_clk _02637_ VGND VGND VPWR VPWR per_uart.uart0.tx_wr sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09092_ _04671_ _04803_ VGND VGND VPWR VPWR _04804_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold900 CPU.registerFile\[22\]\[19\] VGND VGND VPWR VPWR net2141 sky130_fd_sc_hd__dlygate4sd3_1
Xhold911 CPU.registerFile\[17\]\[0\] VGND VGND VPWR VPWR net2152 sky130_fd_sc_hd__dlygate4sd3_1
Xhold922 CPU.registerFile\[31\]\[16\] VGND VGND VPWR VPWR net2163 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold933 CPU.registerFile\[11\]\[25\] VGND VGND VPWR VPWR net2174 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold944 CPU.registerFile\[18\]\[28\] VGND VGND VPWR VPWR net2185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold955 CPU.registerFile\[24\]\[0\] VGND VGND VPWR VPWR net2196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 CPU.registerFile\[16\]\[24\] VGND VGND VPWR VPWR net2207 sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 CPU.registerFile\[24\]\[17\] VGND VGND VPWR VPWR net2218 sky130_fd_sc_hd__dlygate4sd3_1
X_09994_ _05549_ net1892 _05581_ VGND VGND VPWR VPWR _05590_ sky130_fd_sc_hd__mux2_1
Xhold988 CPU.registerFile\[19\]\[21\] VGND VGND VPWR VPWR net2229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold999 CPU.registerFile\[8\]\[21\] VGND VGND VPWR VPWR net2240 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__08368_ _08368_ VGND VGND VPWR VPWR clknet_0__08368_ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_4_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08945_ CPU.Bimm\[4\] VGND VGND VPWR VPWR _04665_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_86_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f__07219_ clknet_0__07219_ VGND VGND VPWR VPWR clknet_1_1__leaf__07219_
+ sky130_fd_sc_hd__clkbuf_16
X_08876_ _04578_ _04595_ VGND VGND VPWR VPWR _04596_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__02721_ clknet_0__02721_ VGND VGND VPWR VPWR clknet_1_0__leaf__02721_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__02652_ clknet_0__02652_ VGND VGND VPWR VPWR clknet_1_0__leaf__02652_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09428_ net2525 _05130_ _04983_ VGND VGND VPWR VPWR _05131_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_23_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_910 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09359_ _05061_ _05052_ _05051_ _05064_ VGND VGND VPWR VPWR _05065_ sky130_fd_sc_hd__or4b_4
XFILLER_0_151_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12370_ _07002_ VGND VGND VPWR VPWR _01401_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11321_ _05514_ net2258 _06371_ VGND VGND VPWR VPWR _06373_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15145__1173 clknet_1_1__leaf__02745_ VGND VGND VPWR VPWR net1205 sky130_fd_sc_hd__inv_2
XFILLER_0_132_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11252_ _06336_ VGND VGND VPWR VPWR _01891_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10203_ _05711_ VGND VGND VPWR VPWR _02330_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11183_ _05511_ net1758 _06299_ VGND VGND VPWR VPWR _06300_ sky130_fd_sc_hd__mux2_1
X_10134_ net1694 _05402_ _05655_ VGND VGND VPWR VPWR _05665_ sky130_fd_sc_hd__mux2_1
X_15991_ _03022_ _03470_ _03471_ _03472_ _02895_ VGND VGND VPWR VPWR _03473_ sky130_fd_sc_hd__o221a_1
X_17730_ net919 _02014_ VGND VGND VPWR VPWR CPU.registerFile\[6\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_10065_ net2010 _05402_ _05618_ VGND VGND VPWR VPWR _05628_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__03968_ clknet_0__03968_ VGND VGND VPWR VPWR clknet_1_0__leaf__03968_
+ sky130_fd_sc_hd__clkbuf_16
X_17661_ net850 _01949_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14873_ clknet_1_1__leaf__02697_ VGND VGND VPWR VPWR _02703_ sky130_fd_sc_hd__buf_1
X_16612_ _03981_ VGND VGND VPWR VPWR _02543_ sky130_fd_sc_hd__clkbuf_1
X_13824_ _07370_ _08238_ VGND VGND VPWR VPWR _08239_ sky130_fd_sc_hd__or2_1
X_17592_ net781 _01880_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10967_ net2098 _05681_ _06179_ VGND VGND VPWR VPWR _06185_ sky130_fd_sc_hd__mux2_1
X_13755_ _07231_ _08169_ _08172_ VGND VGND VPWR VPWR _08173_ sky130_fd_sc_hd__or3_1
Xclkbuf_1_0__f__08357_ clknet_0__08357_ VGND VGND VPWR VPWR clknet_1_0__leaf__08357_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_156_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12706_ net1348 _07187_ VGND VGND VPWR VPWR _07188_ sky130_fd_sc_hd__or2_1
XFILLER_0_155_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16474_ _03252_ _03933_ _03941_ _02935_ VGND VGND VPWR VPWR _03942_ sky130_fd_sc_hd__o211a_1
XFILLER_0_155_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10898_ _06148_ VGND VGND VPWR VPWR _02057_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13686_ CPU.registerFile\[15\]\[23\] _07403_ _07404_ CPU.registerFile\[11\]\[23\]
+ _07405_ VGND VGND VPWR VPWR _08106_ sky130_fd_sc_hd__o221a_1
XFILLER_0_85_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18213_ net54 _02493_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15425_ _02858_ _02919_ _02921_ _08397_ VGND VGND VPWR VPWR _02922_ sky130_fd_sc_hd__a211o_1
XFILLER_0_155_466 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14321__462 clknet_1_1__leaf__08465_ VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__inv_2
XFILLER_0_72_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12637_ net1525 _07142_ VGND VGND VPWR VPWR _00044_ sky130_fd_sc_hd__xor2_1
XFILLER_0_143_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18144_ clknet_leaf_27_clk _02424_ VGND VGND VPWR VPWR CPU.aluIn1\[10\] sky130_fd_sc_hd__dfxtp_2
X_12568_ _07084_ VGND VGND VPWR VPWR _07107_ sky130_fd_sc_hd__buf_4
X_15356_ _05069_ VGND VGND VPWR VPWR _02854_ sky130_fd_sc_hd__buf_4
XFILLER_0_41_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_152_Right_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14307_ clknet_1_1__leaf__08433_ VGND VGND VPWR VPWR _08464_ sky130_fd_sc_hd__buf_1
XFILLER_0_25_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11519_ _06481_ VGND VGND VPWR VPWR _01765_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18075_ net138 _02355_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12499_ _07070_ VGND VGND VPWR VPWR _01340_ sky130_fd_sc_hd__clkbuf_1
X_15287_ _02758_ VGND VGND VPWR VPWR _02786_ sky130_fd_sc_hd__buf_4
Xhold207 mapped_spi_ram.rcv_data\[21\] VGND VGND VPWR VPWR net1448 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold218 mapped_spi_flash.snd_bitcount\[2\] VGND VGND VPWR VPWR net1459 sky130_fd_sc_hd__dlygate4sd3_1
X_17026_ net284 _01348_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[20\] sky130_fd_sc_hd__dfxtp_1
Xhold229 mapped_spi_flash.rcv_data\[1\] VGND VGND VPWR VPWR net1470 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__02715_ _02715_ VGND VGND VPWR VPWR clknet_0__02715_ sky130_fd_sc_hd__clkbuf_16
X_14169_ CPU.Bimm\[7\] _08421_ _08413_ VGND VGND VPWR VPWR _08422_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08730_ _04245_ _04244_ VGND VGND VPWR VPWR _04450_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_147_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17928_ net1117 _02212_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[8\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_0_Left_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08661_ CPU.aluIn1\[23\] VGND VGND VPWR VPWR _04381_ sky130_fd_sc_hd__inv_2
X_17859_ net1048 _02143_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_12762__212 clknet_1_1__leaf__07224_ VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__inv_2
X_08592_ _04310_ _04283_ _04311_ VGND VGND VPWR VPWR _04312_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_85_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14404__537 clknet_1_1__leaf__02656_ VGND VGND VPWR VPWR net569 sky130_fd_sc_hd__inv_2
XFILLER_0_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09213_ CPU.PC\[16\] CPU.PC\[15\] _04924_ VGND VGND VPWR VPWR _04925_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_133_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09144_ _04854_ _04855_ VGND VGND VPWR VPWR _04856_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09075_ _04350_ _04787_ VGND VGND VPWR VPWR _04788_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_114_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold730 CPU.registerFile\[27\]\[11\] VGND VGND VPWR VPWR net1971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 CPU.registerFile\[1\]\[27\] VGND VGND VPWR VPWR net1982 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold752 CPU.registerFile\[27\]\[10\] VGND VGND VPWR VPWR net1993 sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 CPU.registerFile\[17\]\[30\] VGND VGND VPWR VPWR net2004 sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 CPU.registerFile\[7\]\[30\] VGND VGND VPWR VPWR net2015 sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 CPU.registerFile\[19\]\[8\] VGND VGND VPWR VPWR net2026 sky130_fd_sc_hd__dlygate4sd3_1
X_14450__579 clknet_1_0__leaf__02660_ VGND VGND VPWR VPWR net611 sky130_fd_sc_hd__inv_2
Xhold796 CPU.registerFile\[17\]\[16\] VGND VGND VPWR VPWR net2037 sky130_fd_sc_hd__dlygate4sd3_1
X_09977_ _05558_ VGND VGND VPWR VPWR _05581_ sky130_fd_sc_hd__clkbuf_4
X_08928_ mapped_spi_ram.rcv_data\[15\] net19 _04618_ mapped_spi_flash.rcv_data\[15\]
+ VGND VGND VPWR VPWR _04648_ sky130_fd_sc_hd__a22oi_4
X_08859_ _04572_ _04575_ VGND VGND VPWR VPWR _04579_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_28_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11870_ CPU.registerFile\[10\]\[9\] _05717_ _06697_ VGND VGND VPWR VPWR _06700_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__02704_ clknet_0__02704_ VGND VGND VPWR VPWR clknet_1_0__leaf__02704_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15061__1127 clknet_1_0__leaf__02722_ VGND VGND VPWR VPWR net1159 sky130_fd_sc_hd__inv_2
X_10821_ _06107_ VGND VGND VPWR VPWR _02093_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13540_ CPU.registerFile\[6\]\[19\] CPU.registerFile\[7\]\[19\] _07371_ VGND VGND
+ VPWR VPWR _07964_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10752_ _05487_ net1918 _06070_ VGND VGND VPWR VPWR _06071_ sky130_fd_sc_hd__mux2_1
X_14379__514 clknet_1_0__leaf__02654_ VGND VGND VPWR VPWR net546 sky130_fd_sc_hd__inv_2
XFILLER_0_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13471_ CPU.registerFile\[30\]\[17\] CPU.registerFile\[26\]\[17\] _04939_ VGND VGND
+ VPWR VPWR _07897_ sky130_fd_sc_hd__mux2_1
X_10683_ _06033_ VGND VGND VPWR VPWR _06034_ sky130_fd_sc_hd__buf_4
XFILLER_0_109_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12422_ _05090_ net2163 _07024_ VGND VGND VPWR VPWR _07030_ sky130_fd_sc_hd__mux2_1
X_16190_ CPU.registerFile\[5\]\[23\] CPU.registerFile\[4\]\[23\] net15 VGND VGND VPWR
+ VPWR _03666_ sky130_fd_sc_hd__mux2_1
X_12353_ _06993_ VGND VGND VPWR VPWR _01409_ sky130_fd_sc_hd__clkbuf_1
X_15141_ clknet_1_0__leaf__02720_ VGND VGND VPWR VPWR _02745_ sky130_fd_sc_hd__buf_1
XFILLER_0_106_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11304_ _05497_ net2199 _06360_ VGND VGND VPWR VPWR _06364_ sky130_fd_sc_hd__mux2_1
X_12284_ _06948_ VGND VGND VPWR VPWR _01433_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11235_ _06327_ VGND VGND VPWR VPWR _01899_ sky130_fd_sc_hd__clkbuf_1
X_14845__934 clknet_1_1__leaf__02700_ VGND VGND VPWR VPWR net966 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_52_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11166_ _05495_ net2335 _06288_ VGND VGND VPWR VPWR _06291_ sky130_fd_sc_hd__mux2_1
X_10117_ _05656_ VGND VGND VPWR VPWR _02361_ sky130_fd_sc_hd__clkbuf_1
X_11097_ _06254_ VGND VGND VPWR VPWR _01964_ sky130_fd_sc_hd__clkbuf_1
X_15974_ _03065_ _03455_ _03456_ VGND VGND VPWR VPWR _03457_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_147_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17713_ net902 _00011_ VGND VGND VPWR VPWR mapped_spi_ram.state\[3\] sky130_fd_sc_hd__dfxtp_1
X_10048_ _05619_ VGND VGND VPWR VPWR _02393_ sky130_fd_sc_hd__clkbuf_1
Xhold90 _01701_ VGND VGND VPWR VPWR net1331 sky130_fd_sc_hd__dlygate4sd3_1
X_17644_ net833 _01932_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13807_ CPU.registerFile\[8\]\[27\] CPU.registerFile\[12\]\[27\] _07339_ VGND VGND
+ VPWR VPWR _08223_ sky130_fd_sc_hd__mux2_1
X_17575_ net764 _01863_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_11999_ _05170_ net1634 _06758_ VGND VGND VPWR VPWR _06768_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13738_ _07801_ _08153_ _08155_ _07305_ VGND VGND VPWR VPWR _08156_ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14891__976 clknet_1_0__leaf__02704_ VGND VGND VPWR VPWR net1008 sky130_fd_sc_hd__inv_2
XFILLER_0_27_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16457_ _02901_ _03920_ _03925_ _02903_ VGND VGND VPWR VPWR _03926_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_80_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13669_ CPU.registerFile\[16\]\[23\] CPU.registerFile\[20\]\[23\] _07315_ VGND VGND
+ VPWR VPWR _08089_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15408_ CPU.aluIn1\[1\] _07705_ _02880_ _02905_ _07737_ VGND VGND VPWR VPWR _02415_
+ sky130_fd_sc_hd__o221a_1
X_16388_ _02827_ _03857_ _03858_ VGND VGND VPWR VPWR _03859_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18127_ net190 _02407_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[25\] sky130_fd_sc_hd__dfxtp_1
X_15339_ _02827_ _02830_ _02837_ VGND VGND VPWR VPWR _02838_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_151_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18058_ net1231 _02338_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17009_ net267 _01331_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_09900_ _05208_ VGND VGND VPWR VPWR _05535_ sky130_fd_sc_hd__buf_4
XFILLER_0_21_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09831_ _04658_ VGND VGND VPWR VPWR _05487_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_111_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09762_ _04660_ _04661_ VGND VGND VPWR VPWR _05450_ sky130_fd_sc_hd__nand2_4
X_08713_ _04432_ VGND VGND VPWR VPWR _04433_ sky130_fd_sc_hd__inv_2
X_09693_ mapped_spi_ram.rcv_data\[10\] _04783_ _04784_ mapped_spi_flash.rcv_data\[10\]
+ VGND VGND VPWR VPWR _05384_ sky130_fd_sc_hd__a22o_4
XFILLER_0_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer11 net1253 VGND VGND VPWR VPWR net1252 sky130_fd_sc_hd__dlygate4sd1_1
X_08644_ _04228_ _04363_ VGND VGND VPWR VPWR _04364_ sky130_fd_sc_hd__or2_4
Xrebuffer22 net1264 VGND VGND VPWR VPWR net1263 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer33 _04542_ VGND VGND VPWR VPWR net1287 sky130_fd_sc_hd__clkbuf_2
Xrebuffer44 net1292 VGND VGND VPWR VPWR net1291 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15144__1172 clknet_1_0__leaf__02745_ VGND VGND VPWR VPWR net1204 sky130_fd_sc_hd__inv_2
X_08575_ CPU.instr\[3\] CPU.instr\[2\] _04292_ net1275 VGND VGND VPWR VPWR _04295_
+ sky130_fd_sc_hd__nor4b_2
XFILLER_0_49_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_876 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_147_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_697 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15229__139 clknet_1_1__leaf__02753_ VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__inv_2
XFILLER_0_44_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09127_ CPU.PC\[17\] _04838_ VGND VGND VPWR VPWR _04839_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_98_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_801 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09058_ _04353_ _04489_ _04771_ VGND VGND VPWR VPWR _04772_ sky130_fd_sc_hd__a21o_1
X_14003__284 clknet_1_0__leaf__08360_ VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__inv_2
XFILLER_0_130_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold560 CPU.registerFile\[14\]\[28\] VGND VGND VPWR VPWR net1801 sky130_fd_sc_hd__dlygate4sd3_1
Xhold571 CPU.registerFile\[19\]\[20\] VGND VGND VPWR VPWR net1812 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ _06212_ VGND VGND VPWR VPWR _01999_ sky130_fd_sc_hd__clkbuf_1
Xhold582 CPU.registerFile\[27\]\[9\] VGND VGND VPWR VPWR net1823 sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 CPU.registerFile\[30\]\[28\] VGND VGND VPWR VPWR net1834 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ _07296_ VGND VGND VPWR VPWR _07412_ sky130_fd_sc_hd__buf_4
Xhold1260 CPU.registerFile\[24\]\[8\] VGND VGND VPWR VPWR net2501 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1271 CPU.registerFile\[25\]\[16\] VGND VGND VPWR VPWR net2512 sky130_fd_sc_hd__dlygate4sd3_1
X_11922_ _06727_ VGND VGND VPWR VPWR _01609_ sky130_fd_sc_hd__clkbuf_1
Xhold1282 CPU.registerFile\[10\]\[0\] VGND VGND VPWR VPWR net2523 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1293 CPU.registerFile\[13\]\[15\] VGND VGND VPWR VPWR net2534 sky130_fd_sc_hd__dlygate4sd3_1
X_15690_ _02818_ _03179_ _03180_ VGND VGND VPWR VPWR _03181_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_400 _07250_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_411 _04659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ CPU.registerFile\[10\]\[17\] _05700_ _06686_ VGND VGND VPWR VPWR _06691_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_157_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17360_ net549 _01648_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_10804_ _05543_ net1746 _06092_ VGND VGND VPWR VPWR _06098_ sky130_fd_sc_hd__mux2_1
X_11784_ _06654_ VGND VGND VPWR VPWR _01674_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16311_ _02796_ _03783_ VGND VGND VPWR VPWR _03784_ sky130_fd_sc_hd__or2_1
X_13523_ _07398_ _07946_ _07947_ VGND VGND VPWR VPWR _07948_ sky130_fd_sc_hd__o21a_1
X_17291_ net480 _01579_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_10735_ _06061_ VGND VGND VPWR VPWR _02133_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_45_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16242_ CPU.registerFile\[6\]\[24\] _03057_ _03140_ _03716_ VGND VGND VPWR VPWR _03717_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_745 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13454_ _07412_ _07879_ _07880_ VGND VGND VPWR VPWR _07881_ sky130_fd_sc_hd__o21a_1
X_10666_ mapped_spi_flash.rcv_bitcount\[4\] _05964_ VGND VGND VPWR VPWR _06023_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12405_ _04798_ net2254 _07013_ VGND VGND VPWR VPWR _07021_ sky130_fd_sc_hd__mux2_1
X_16173_ _03252_ _03640_ _03649_ _08408_ VGND VGND VPWR VPWR _03650_ sky130_fd_sc_hd__o211a_1
X_13385_ CPU.registerFile\[21\]\[14\] _07244_ _07429_ CPU.registerFile\[17\]\[14\]
+ _07349_ VGND VGND VPWR VPWR _07814_ sky130_fd_sc_hd__o221a_1
X_10597_ net1443 _05968_ _05979_ _05980_ VGND VGND VPWR VPWR _02189_ sky130_fd_sc_hd__o211a_1
X_12336_ _06984_ VGND VGND VPWR VPWR _01417_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12267_ _06935_ VGND VGND VPWR VPWR _01437_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14433__563 clknet_1_1__leaf__02659_ VGND VGND VPWR VPWR net595 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_149_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11218_ _05547_ net1989 _06310_ VGND VGND VPWR VPWR _06318_ sky130_fd_sc_hd__mux2_1
X_12198_ _06882_ VGND VGND VPWR VPWR _01453_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11149_ _06281_ VGND VGND VPWR VPWR _01939_ sky130_fd_sc_hd__clkbuf_1
X_15957_ CPU.registerFile\[30\]\[16\] CPU.registerFile\[26\]\[16\] _03247_ VGND VGND
+ VPWR VPWR _03440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_618 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15888_ _02771_ _03370_ _03371_ _03372_ _02807_ VGND VGND VPWR VPWR _03373_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_90_Left_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17627_ net816 _01915_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[13\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_82_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17558_ net747 _01846_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15019__1091 clknet_1_1__leaf__02717_ VGND VGND VPWR VPWR net1123 sky130_fd_sc_hd__inv_2
XFILLER_0_73_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17489_ net678 _01777_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_16585__57 clknet_1_1__leaf__03969_ VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__inv_2
XFILLER_0_129_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14516__638 clknet_1_0__leaf__02667_ VGND VGND VPWR VPWR net670 sky130_fd_sc_hd__inv_2
XFILLER_0_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14254__426 clknet_1_0__leaf__08435_ VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__inv_2
X_15060__1126 clknet_1_0__leaf__02722_ VGND VGND VPWR VPWR net1158 sky130_fd_sc_hd__inv_2
XFILLER_0_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09814_ _05478_ VGND VGND VPWR VPWR _02518_ sky130_fd_sc_hd__clkbuf_1
X_09745_ _04504_ _04208_ _05433_ VGND VGND VPWR VPWR _05434_ sky130_fd_sc_hd__nand3_1
XPHY_EDGE_ROW_129_Left_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09676_ _04289_ _04304_ _04306_ VGND VGND VPWR VPWR _05368_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08627_ _04346_ _04244_ _04242_ _04240_ VGND VGND VPWR VPWR _04347_ sky130_fd_sc_hd__a31o_4
XTAP_TAPCELL_ROW_124_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08558_ _04277_ VGND VGND VPWR VPWR _04278_ sky130_fd_sc_hd__inv_2
X_14874__960 clknet_1_1__leaf__02703_ VGND VGND VPWR VPWR net992 sky130_fd_sc_hd__inv_2
XFILLER_0_92_610 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08489_ _04208_ CPU.Jimm\[14\] CPU.Jimm\[13\] VGND VGND VPWR VPWR _04209_ sky130_fd_sc_hd__and3b_1
XFILLER_0_92_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10520_ net1354 _05887_ _05856_ _05924_ VGND VGND VPWR VPWR _05925_ sky130_fd_sc_hd__a211o_1
XFILLER_0_80_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_138_Left_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10451_ net1399 _05850_ _05851_ _05865_ VGND VGND VPWR VPWR _05866_ sky130_fd_sc_hd__a211o_1
XFILLER_0_122_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13170_ CPU.registerFile\[16\]\[8\] CPU.registerFile\[20\]\[8\] _07233_ VGND VGND
+ VPWR VPWR _07605_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10382_ net2540 VGND VGND VPWR VPWR _05814_ sky130_fd_sc_hd__inv_2
X_12121_ _05027_ net2442 _06830_ VGND VGND VPWR VPWR _06833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12052_ _06796_ VGND VGND VPWR VPWR _01547_ sky130_fd_sc_hd__clkbuf_1
Xhold390 CPU.registerFile\[18\]\[19\] VGND VGND VPWR VPWR net1631 sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ net1583 _05717_ _06201_ VGND VGND VPWR VPWR _06204_ sky130_fd_sc_hd__mux2_1
X_16860_ _04148_ per_uart.rx_error _04137_ _03975_ VGND VGND VPWR VPWR _04149_ sky130_fd_sc_hd__a22o_1
X_15811_ CPU.aluIn1\[11\] _03081_ _03298_ _03080_ VGND VGND VPWR VPWR _02425_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_144_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_144_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16791_ _05288_ _08454_ _04952_ VGND VGND VPWR VPWR _04102_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15742_ CPU.registerFile\[2\]\[10\] _03227_ _03228_ CPU.registerFile\[3\]\[10\] _03230_
+ VGND VGND VPWR VPWR _03231_ sky130_fd_sc_hd__a221o_1
X_12954_ _07394_ VGND VGND VPWR VPWR _07395_ sky130_fd_sc_hd__buf_2
Xhold1090 CPU.registerFile\[19\]\[24\] VGND VGND VPWR VPWR net2331 sky130_fd_sc_hd__dlygate4sd3_1
X_11905_ _06718_ VGND VGND VPWR VPWR _01617_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15673_ CPU.registerFile\[13\]\[8\] _03123_ VGND VGND VPWR VPWR _03164_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_47_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ _05308_ VGND VGND VPWR VPWR _07327_ sky130_fd_sc_hd__clkbuf_8
XANTENNA_230 clknet_1_1__leaf__02693_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_241 _03021_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_252 _05026_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17412_ net601 _01700_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[5\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_263 _05129_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_114_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11836_ net2273 _05683_ _06675_ VGND VGND VPWR VPWR _06682_ sky130_fd_sc_hd__mux2_1
XANTENNA_274 _05543_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_285 _05594_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_296 _07271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17343_ net532 _01631_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11767_ _06645_ VGND VGND VPWR VPWR _01682_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_60_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13506_ CPU.registerFile\[5\]\[18\] CPU.registerFile\[4\]\[18\] _07577_ VGND VGND
+ VPWR VPWR _07931_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17274_ net463 _01562_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_10718_ _06052_ VGND VGND VPWR VPWR _02141_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11698_ mapped_spi_ram.rcv_data\[11\] _06590_ _06602_ _06594_ VGND VGND VPWR VPWR
+ _01707_ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16225_ CPU.registerFile\[8\]\[24\] _02789_ _03117_ _03699_ VGND VGND VPWR VPWR _03700_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13437_ CPU.registerFile\[18\]\[16\] CPU.registerFile\[22\]\[16\] _07258_ VGND VGND
+ VPWR VPWR _07864_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_155_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer2 net1246 VGND VGND VPWR VPWR net1243 sky130_fd_sc_hd__clkbuf_2
X_10649_ net3 _05967_ _06009_ _06006_ VGND VGND VPWR VPWR _02166_ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_140_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16156_ CPU.registerFile\[14\]\[22\] CPU.registerFile\[10\]\[22\] _02906_ VGND VGND
+ VPWR VPWR _03633_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13368_ _07570_ _07794_ _07795_ _07797_ _04814_ VGND VGND VPWR VPWR _07798_ sky130_fd_sc_hd__a221o_1
X_15107_ _07192_ _02740_ _02726_ VGND VGND VPWR VPWR _02283_ sky130_fd_sc_hd__a21oi_1
X_12319_ net2270 _06974_ _06861_ VGND VGND VPWR VPWR _06975_ sky130_fd_sc_hd__mux2_1
X_15143__1171 clknet_1_1__leaf__02745_ VGND VGND VPWR VPWR net1203 sky130_fd_sc_hd__inv_2
X_16087_ CPU.registerFile\[1\]\[20\] _03228_ _03565_ _02818_ VGND VGND VPWR VPWR _03566_
+ sky130_fd_sc_hd__a22o_1
X_13299_ _07398_ _07729_ _07730_ VGND VGND VPWR VPWR _07731_ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15038_ _07123_ _04193_ _04492_ VGND VGND VPWR VPWR _02719_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_75_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14704__808 clknet_1_0__leaf__02685_ VGND VGND VPWR VPWR net840 sky130_fd_sc_hd__inv_2
X_16989_ clknet_leaf_21_clk _01315_ VGND VGND VPWR VPWR CPU.rs2\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09530_ _04974_ _05225_ _05226_ _04955_ _05227_ VGND VGND VPWR VPWR _05228_ sky130_fd_sc_hd__o221a_1
X_09461_ _05158_ _05161_ _04373_ VGND VGND VPWR VPWR _05162_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_35_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09392_ CPU.PC\[15\] _04924_ VGND VGND VPWR VPWR _05096_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_789 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_681 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09728_ _05415_ _05417_ VGND VGND VPWR VPWR _05418_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09659_ _04287_ _04307_ VGND VGND VPWR VPWR _05352_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12670_ net1433 _07160_ VGND VGND VPWR VPWR _07163_ sky130_fd_sc_hd__nor2_1
X_16549__24 clknet_1_1__leaf__03966_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__inv_2
XFILLER_0_65_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11621_ mapped_spi_ram.snd_bitcount\[4\] _06550_ VGND VGND VPWR VPWR _06551_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_146_Left_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14340_ clknet_1_0__leaf__08433_ VGND VGND VPWR VPWR _08467_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_42_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11552_ _06501_ _05872_ VGND VGND VPWR VPWR _06504_ sky130_fd_sc_hd__nor2_1
X_16564__38 clknet_1_1__leaf__03967_ VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10503_ _04516_ net1243 _04515_ _04629_ VGND VGND VPWR VPWR _05910_ sky130_fd_sc_hd__a31o_1
X_14271_ _04483_ _04218_ VGND VGND VPWR VPWR _08450_ sky130_fd_sc_hd__nand2_1
X_11483_ _05539_ net2429 _06455_ VGND VGND VPWR VPWR _06459_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16010_ CPU.registerFile\[28\]\[17\] CPU.registerFile\[24\]\[17\] _02918_ VGND VGND
+ VPWR VPWR _03492_ sky130_fd_sc_hd__mux2_1
X_10434_ net1374 _05850_ _05851_ _05853_ VGND VGND VPWR VPWR _05854_ sky130_fd_sc_hd__a211o_1
X_13222_ _07653_ _07654_ _07655_ VGND VGND VPWR VPWR _07656_ sky130_fd_sc_hd__o21ai_2
X_14237__410 clknet_1_0__leaf__08434_ VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__inv_2
XFILLER_0_60_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10365_ _05804_ VGND VGND VPWR VPWR _02246_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13153_ _07475_ _07587_ _07588_ VGND VGND VPWR VPWR _07589_ sky130_fd_sc_hd__o21a_1
XFILLER_0_150_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12104_ _04748_ net2292 _06819_ VGND VGND VPWR VPWR _06824_ sky130_fd_sc_hd__mux2_1
X_17961_ net1149 _02245_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_13084_ CPU.registerFile\[13\]\[5\] _07281_ _07521_ CPU.registerFile\[9\]\[5\] _07285_
+ VGND VGND VPWR VPWR _07522_ sky130_fd_sc_hd__o221a_1
X_10296_ _05767_ VGND VGND VPWR VPWR _02293_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_155_Left_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12035_ _06787_ VGND VGND VPWR VPWR _01555_ sky130_fd_sc_hd__clkbuf_1
X_16912_ net1750 _04182_ VGND VGND VPWR VPWR _04185_ sky130_fd_sc_hd__or2_1
X_17892_ net1081 _02176_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[10\] sky130_fd_sc_hd__dfxtp_1
X_15018__1090 clknet_1_0__leaf__02717_ VGND VGND VPWR VPWR net1122 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16843_ net1508 per_uart.rx_data\[0\] _04139_ VGND VGND VPWR VPWR _04140_ sky130_fd_sc_hd__mux2_1
X_14545__664 clknet_1_0__leaf__02670_ VGND VGND VPWR VPWR net696 sky130_fd_sc_hd__inv_2
X_16774_ _04052_ _05024_ _08453_ VGND VGND VPWR VPWR _04088_ sky130_fd_sc_hd__or3b_1
XFILLER_0_88_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15725_ _02848_ _03210_ _03214_ _02843_ VGND VGND VPWR VPWR _03215_ sky130_fd_sc_hd__a211o_1
XFILLER_0_158_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12937_ _07369_ _07372_ _07377_ _07231_ VGND VGND VPWR VPWR _07378_ sky130_fd_sc_hd__a211o_4
XFILLER_0_76_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15656_ CPU.registerFile\[1\]\[7\] _02814_ _03147_ _02943_ VGND VGND VPWR VPWR _03148_
+ sky130_fd_sc_hd__a22o_1
X_12868_ CPU.mem_wdata\[0\] _07229_ _07310_ _07135_ VGND VGND VPWR VPWR _01295_ sky130_fd_sc_hd__o211a_1
XFILLER_0_158_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14607_ clknet_1_1__leaf__02675_ VGND VGND VPWR VPWR _02677_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_157_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11819_ _06672_ VGND VGND VPWR VPWR _01657_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_157_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15587_ CPU.aluIn1\[5\] _08018_ _03079_ _03080_ VGND VGND VPWR VPWR _02419_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12799_ _05338_ _07241_ VGND VGND VPWR VPWR _07242_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17326_ net515 _01614_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_126_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f__03964_ clknet_0__03964_ VGND VGND VPWR VPWR clknet_1_1__leaf__03964_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_83_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17257_ net447 _01545_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[18\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_77_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16208_ CPU.registerFile\[15\]\[23\] CPU.registerFile\[11\]\[23\] _03247_ VGND VGND
+ VPWR VPWR _03684_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17188_ clknet_leaf_26_clk _01476_ VGND VGND VPWR VPWR CPU.Jimm\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14710__812 clknet_1_0__leaf__02687_ VGND VGND VPWR VPWR net844 sky130_fd_sc_hd__inv_2
X_16139_ CPU.registerFile\[7\]\[21\] _03317_ VGND VGND VPWR VPWR _03617_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14290__434 clknet_1_1__leaf__08462_ VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__inv_2
XFILLER_0_110_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08961_ _04672_ _04674_ _04676_ _04679_ VGND VGND VPWR VPWR _04680_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_90_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14628__739 clknet_1_0__leaf__02678_ VGND VGND VPWR VPWR net771 sky130_fd_sc_hd__inv_2
X_08892_ _04608_ _04611_ VGND VGND VPWR VPWR _04612_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_108_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09513_ mapped_spi_flash.rcv_data\[17\] _04709_ _04644_ per_uart.tx_busy VGND VGND
+ VPWR VPWR _05211_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_88_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09444_ _05143_ _05145_ _04374_ VGND VGND VPWR VPWR _05146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09375_ _04441_ _05079_ VGND VGND VPWR VPWR _05080_ sky130_fd_sc_hd__and2b_1
XFILLER_0_148_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10150_ net1842 _05675_ _05671_ VGND VGND VPWR VPWR _05676_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10081_ _05637_ VGND VGND VPWR VPWR _02378_ sky130_fd_sc_hd__clkbuf_1
X_13840_ _07650_ _08253_ _08254_ VGND VGND VPWR VPWR _08255_ sky130_fd_sc_hd__o21ai_1
X_13771_ _08184_ _08187_ _07584_ VGND VGND VPWR VPWR _08188_ sky130_fd_sc_hd__a21oi_2
X_10983_ _06193_ VGND VGND VPWR VPWR _02017_ sky130_fd_sc_hd__clkbuf_1
X_15510_ CPU.registerFile\[5\]\[4\] CPU.registerFile\[4\]\[4\] _02806_ VGND VGND VPWR
+ VPWR _03005_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12722_ per_uart.d_in_uart\[6\] _07178_ _07203_ net1410 VGND VGND VPWR VPWR _07204_
+ sky130_fd_sc_hd__a22o_1
X_16490_ CPU.registerFile\[30\]\[31\] _05050_ _02770_ _03957_ VGND VGND VPWR VPWR
+ _03958_ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15142__1170 clknet_1_0__leaf__02745_ VGND VGND VPWR VPWR net1202 sky130_fd_sc_hd__inv_2
XFILLER_0_139_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15441_ CPU.registerFile\[6\]\[2\] _02870_ _02894_ _02937_ VGND VGND VPWR VPWR _02938_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_127_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_133_Right_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12653_ CPU.cycles\[13\] _07150_ net1487 VGND VGND VPWR VPWR _07153_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_139_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18160_ clknet_leaf_29_clk _02440_ VGND VGND VPWR VPWR CPU.aluIn1\[26\] sky130_fd_sc_hd__dfxtp_2
X_11604_ net1388 _06501_ _06496_ CPU.mem_wdata\[6\] _06508_ VGND VGND VPWR VPWR _06541_
+ sky130_fd_sc_hd__a221o_1
X_15372_ _08395_ VGND VGND VPWR VPWR _02870_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_136_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12584_ _07115_ VGND VGND VPWR VPWR _01267_ sky130_fd_sc_hd__clkbuf_1
X_17111_ clknet_leaf_23_clk _00044_ VGND VGND VPWR VPWR CPU.cycles\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_646 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18091_ net154 _02371_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_11535_ _05816_ net1313 _06489_ _06492_ net1319 VGND VGND VPWR VPWR _01760_ sky130_fd_sc_hd__a32o_1
XFILLER_0_135_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_819 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__02700_ clknet_0__02700_ VGND VGND VPWR VPWR clknet_1_1__leaf__02700_
+ sky130_fd_sc_hd__clkbuf_16
X_17042_ net300 _01364_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_152_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_152_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11466_ _05522_ net2512 _06444_ VGND VGND VPWR VPWR _06450_ sky130_fd_sc_hd__mux2_1
X_13205_ _07638_ VGND VGND VPWR VPWR _07639_ sky130_fd_sc_hd__clkbuf_4
X_10417_ _05825_ VGND VGND VPWR VPWR _05841_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11397_ _06413_ VGND VGND VPWR VPWR _01823_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__02662_ _02662_ VGND VGND VPWR VPWR clknet_0__02662_ sky130_fd_sc_hd__clkbuf_16
X_13136_ _07245_ _07571_ VGND VGND VPWR VPWR _07572_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_55_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10348_ _05795_ VGND VGND VPWR VPWR _02254_ sky130_fd_sc_hd__clkbuf_1
X_10279_ _05758_ VGND VGND VPWR VPWR _02301_ sky130_fd_sc_hd__clkbuf_1
X_17944_ net1133 _02228_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[24\] sky130_fd_sc_hd__dfxtp_1
X_13067_ CPU.registerFile\[16\]\[5\] CPU.registerFile\[20\]\[5\] _07314_ VGND VGND
+ VPWR VPWR _07505_ sky130_fd_sc_hd__mux2_1
X_12018_ _05381_ net1959 _06769_ VGND VGND VPWR VPWR _06778_ sky130_fd_sc_hd__mux2_1
X_17875_ net1064 _02159_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_bitcount\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16826_ _04127_ VGND VGND VPWR VPWR _02611_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16757_ _03995_ _05078_ _07132_ VGND VGND VPWR VPWR _04074_ sky130_fd_sc_hd__o21ai_1
X_15708_ CPU.registerFile\[15\]\[9\] _02826_ _02770_ _03197_ VGND VGND VPWR VPWR _03198_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_598 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16688_ _04010_ _04014_ _04015_ VGND VGND VPWR VPWR _02585_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14816__909 clknet_1_0__leaf__02696_ VGND VGND VPWR VPWR net941 sky130_fd_sc_hd__inv_2
X_14209__386 clknet_1_0__leaf__08430_ VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15639_ CPU.registerFile\[28\]\[7\] _02791_ VGND VGND VPWR VPWR _03131_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09160_ _04499_ CPU.Iimm\[1\] _04660_ _04830_ VGND VGND VPWR VPWR _04872_ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18358_ clknet_leaf_4_clk _02636_ VGND VGND VPWR VPWR per_uart.uart_ctrl\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17309_ net498 _01597_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09091_ _04347_ _04461_ VGND VGND VPWR VPWR _04803_ sky130_fd_sc_hd__xor2_2
X_12756__209 clknet_1_1__leaf__07221_ VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__inv_2
X_18289_ net122 _02569_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16543__19 clknet_1_0__leaf__03965_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__inv_2
XFILLER_0_114_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold901 CPU.registerFile\[1\]\[23\] VGND VGND VPWR VPWR net2142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold912 CPU.registerFile\[29\]\[1\] VGND VGND VPWR VPWR net2153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 CPU.registerFile\[23\]\[29\] VGND VGND VPWR VPWR net2164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold934 CPU.registerFile\[13\]\[8\] VGND VGND VPWR VPWR net2175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold945 CPU.registerFile\[14\]\[9\] VGND VGND VPWR VPWR net2186 sky130_fd_sc_hd__dlygate4sd3_1
Xhold956 CPU.registerFile\[11\]\[7\] VGND VGND VPWR VPWR net2197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 CPU.registerFile\[1\]\[0\] VGND VGND VPWR VPWR net2208 sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 CPU.registerFile\[1\]\[15\] VGND VGND VPWR VPWR net2219 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_896 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold989 CPU.registerFile\[3\]\[28\] VGND VGND VPWR VPWR net2230 sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ _05589_ VGND VGND VPWR VPWR _02450_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__08367_ _08367_ VGND VGND VPWR VPWR clknet_0__08367_ sky130_fd_sc_hd__clkbuf_16
X_08944_ CPU.Bimm\[2\] VGND VGND VPWR VPWR _04664_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_4_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08875_ CPU.aluIn1\[22\] _04496_ VGND VGND VPWR VPWR _04595_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0__f__02720_ clknet_0__02720_ VGND VGND VPWR VPWR clknet_1_0__leaf__02720_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09427_ _05129_ VGND VGND VPWR VPWR _05130_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_23_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09358_ _04916_ _04926_ _05062_ _05063_ _04974_ VGND VGND VPWR VPWR _05064_ sky130_fd_sc_hd__o32a_1
XFILLER_0_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09289_ _04995_ _04997_ _04374_ VGND VGND VPWR VPWR _04998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14574__690 clknet_1_0__leaf__02673_ VGND VGND VPWR VPWR net722 sky130_fd_sc_hd__inv_2
X_11320_ _06372_ VGND VGND VPWR VPWR _01859_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_134_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11251_ CPU.registerFile\[9\]\[21\] _05691_ _06335_ VGND VGND VPWR VPWR _06336_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10202_ net2492 _05710_ _05692_ VGND VGND VPWR VPWR _05711_ sky130_fd_sc_hd__mux2_1
X_11182_ _06287_ VGND VGND VPWR VPWR _06299_ sky130_fd_sc_hd__buf_4
X_10133_ _05664_ VGND VGND VPWR VPWR _02353_ sky130_fd_sc_hd__clkbuf_1
X_15990_ CPU.registerFile\[20\]\[17\] _02855_ _03026_ VGND VGND VPWR VPWR _03472_
+ sky130_fd_sc_hd__a21o_1
X_10064_ _05627_ VGND VGND VPWR VPWR _02385_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__03967_ clknet_0__03967_ VGND VGND VPWR VPWR clknet_1_0__leaf__03967_
+ sky130_fd_sc_hd__clkbuf_16
X_17660_ net849 _01948_ VGND VGND VPWR VPWR CPU.registerFile\[8\]\[14\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_50_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16611_ net2069 net1540 _03979_ VGND VGND VPWR VPWR _03981_ sky130_fd_sc_hd__mux2_1
X_13823_ CPU.registerFile\[14\]\[28\] CPU.registerFile\[10\]\[28\] _04936_ VGND VGND
+ VPWR VPWR _08238_ sky130_fd_sc_hd__mux2_1
X_17591_ net780 _01879_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13754_ _07576_ _08170_ _08171_ _08082_ VGND VGND VPWR VPWR _08172_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10966_ _06184_ VGND VGND VPWR VPWR _02025_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0__f__08356_ clknet_0__08356_ VGND VGND VPWR VPWR clknet_1_0__leaf__08356_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12705_ net1440 _07186_ VGND VGND VPWR VPWR _07187_ sky130_fd_sc_hd__or2_1
X_16473_ _02949_ _03937_ _03940_ VGND VGND VPWR VPWR _03941_ sky130_fd_sc_hd__or3_2
X_13685_ _07398_ _08104_ VGND VGND VPWR VPWR _08105_ sky130_fd_sc_hd__or2_1
X_10897_ net1711 _05679_ _06143_ VGND VGND VPWR VPWR _06148_ sky130_fd_sc_hd__mux2_1
X_18212_ net53 _02492_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15424_ CPU.registerFile\[24\]\[2\] _02816_ _05071_ _02920_ VGND VGND VPWR VPWR _02921_
+ sky130_fd_sc_hd__o211a_1
X_14657__765 clknet_1_0__leaf__02681_ VGND VGND VPWR VPWR net797 sky130_fd_sc_hd__inv_2
XFILLER_0_54_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12636_ _07142_ _07143_ VGND VGND VPWR VPWR _00043_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_478 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18143_ clknet_leaf_27_clk _02423_ VGND VGND VPWR VPWR CPU.aluIn1\[9\] sky130_fd_sc_hd__dfxtp_4
X_15355_ CPU.registerFile\[9\]\[1\] CPU.registerFile\[13\]\[1\] _02852_ VGND VGND
+ VPWR VPWR _02853_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12567_ _07106_ VGND VGND VPWR VPWR _01275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_640 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_124_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18074_ net137 _02354_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_11518_ mapped_spi_flash.div_counter\[0\] _06031_ _04193_ VGND VGND VPWR VPWR _06481_
+ sky130_fd_sc_hd__and3b_1
X_15286_ _02768_ _02783_ _02784_ VGND VGND VPWR VPWR _02785_ sky130_fd_sc_hd__a21o_1
X_12498_ net1827 _05710_ _07060_ VGND VGND VPWR VPWR _07070_ sky130_fd_sc_hd__mux2_1
Xhold208 _01717_ VGND VGND VPWR VPWR net1449 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17025_ net283 _01347_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold219 mapped_spi_ram.rcv_data\[27\] VGND VGND VPWR VPWR net1460 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11449_ _05505_ net2166 _06433_ VGND VGND VPWR VPWR _06441_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__02714_ _02714_ VGND VGND VPWR VPWR clknet_0__02714_ sky130_fd_sc_hd__clkbuf_16
X_14168_ _04744_ VGND VGND VPWR VPWR _08421_ sky130_fd_sc_hd__inv_2
X_13119_ _07235_ VGND VGND VPWR VPWR _07556_ sky130_fd_sc_hd__buf_4
X_14099_ _08377_ VGND VGND VPWR VPWR _01459_ sky130_fd_sc_hd__clkbuf_1
X_17927_ net1116 _02211_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[7\] sky130_fd_sc_hd__dfxtp_1
X_14822__913 clknet_1_0__leaf__02698_ VGND VGND VPWR VPWR net945 sky130_fd_sc_hd__inv_2
X_08660_ _04379_ _04227_ VGND VGND VPWR VPWR _04380_ sky130_fd_sc_hd__nor2_1
X_17858_ net1047 _02142_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_16809_ _06482_ _07198_ _04114_ _04115_ VGND VGND VPWR VPWR _02606_ sky130_fd_sc_hd__a31o_1
X_08591_ _04280_ VGND VGND VPWR VPWR _04311_ sky130_fd_sc_hd__inv_2
X_17789_ net978 _02073_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_85_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09212_ CPU.PC\[14\] _04923_ VGND VGND VPWR VPWR _04924_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09143_ CPU.PC\[11\] _04853_ VGND VGND VPWR VPWR _04855_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09074_ _04382_ _04462_ VGND VGND VPWR VPWR _04787_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_936 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold720 CPU.registerFile\[22\]\[8\] VGND VGND VPWR VPWR net1961 sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 CPU.PC\[13\] VGND VGND VPWR VPWR net1972 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold742 CPU.registerFile\[17\]\[3\] VGND VGND VPWR VPWR net1983 sky130_fd_sc_hd__dlygate4sd3_1
Xhold753 CPU.registerFile\[13\]\[20\] VGND VGND VPWR VPWR net1994 sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 CPU.registerFile\[27\]\[24\] VGND VGND VPWR VPWR net2005 sky130_fd_sc_hd__dlygate4sd3_1
Xhold775 CPU.registerFile\[31\]\[30\] VGND VGND VPWR VPWR net2016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 CPU.registerFile\[20\]\[1\] VGND VGND VPWR VPWR net2027 sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 CPU.registerFile\[18\]\[8\] VGND VGND VPWR VPWR net2038 sky130_fd_sc_hd__dlygate4sd3_1
X_09976_ _05580_ VGND VGND VPWR VPWR _02458_ sky130_fd_sc_hd__clkbuf_1
X_08927_ per_uart.rx_data\[7\] _04643_ _04644_ per_uart.rx_error _04646_ VGND VGND
+ VPWR VPWR _04647_ sky130_fd_sc_hd__a221oi_4
XPHY_EDGE_ROW_110_Left_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08858_ _04576_ _04575_ _04577_ _04572_ VGND VGND VPWR VPWR _04578_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_28_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__02703_ clknet_0__02703_ VGND VGND VPWR VPWR clknet_1_0__leaf__02703_
+ sky130_fd_sc_hd__clkbuf_16
X_08789_ _04507_ _04508_ VGND VGND VPWR VPWR _04509_ sky130_fd_sc_hd__nand2_1
X_10820_ net1598 _05668_ _06106_ VGND VGND VPWR VPWR _06107_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10751_ _06069_ VGND VGND VPWR VPWR _06070_ sky130_fd_sc_hd__buf_4
XFILLER_0_48_782 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13470_ _07653_ _07894_ _07895_ VGND VGND VPWR VPWR _07896_ sky130_fd_sc_hd__o21a_1
X_10682_ _05737_ _06032_ VGND VGND VPWR VPWR _06033_ sky130_fd_sc_hd__nand2_2
X_12421_ _07029_ VGND VGND VPWR VPWR _01377_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12352_ net1244 net2123 _06988_ VGND VGND VPWR VPWR _06993_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11303_ _06363_ VGND VGND VPWR VPWR _01867_ sky130_fd_sc_hd__clkbuf_1
X_15206__118 clknet_1_1__leaf__02751_ VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__inv_2
X_12283_ CPU.aluReg\[9\] _06947_ _06924_ VGND VGND VPWR VPWR _06948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11234_ net2391 _05675_ _06324_ VGND VGND VPWR VPWR _06327_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11165_ _06290_ VGND VGND VPWR VPWR _01932_ sky130_fd_sc_hd__clkbuf_1
X_10116_ net2376 _05188_ _05655_ VGND VGND VPWR VPWR _05656_ sky130_fd_sc_hd__mux2_1
X_11096_ net1582 _05673_ _06252_ VGND VGND VPWR VPWR _06254_ sky130_fd_sc_hd__mux2_1
X_15973_ CPU.registerFile\[16\]\[16\] _02831_ _02834_ CPU.registerFile\[17\]\[16\]
+ _02854_ VGND VGND VPWR VPWR _03456_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_147_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17712_ net901 _00010_ VGND VGND VPWR VPWR mapped_spi_ram.state\[2\] sky130_fd_sc_hd__dfxtp_2
X_10047_ net1966 _05188_ _05618_ VGND VGND VPWR VPWR _05619_ sky130_fd_sc_hd__mux2_1
Xhold80 mapped_spi_ram.cmd_addr\[28\] VGND VGND VPWR VPWR net1321 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 net8 VGND VGND VPWR VPWR net1332 sky130_fd_sc_hd__dlygate4sd3_1
X_17643_ net832 _01931_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13806_ _07818_ _08220_ _08221_ VGND VGND VPWR VPWR _08222_ sky130_fd_sc_hd__o21a_1
XFILLER_0_86_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17574_ net763 _01862_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_11998_ _06767_ VGND VGND VPWR VPWR _01573_ sky130_fd_sc_hd__clkbuf_1
X_13737_ _07987_ _08154_ VGND VGND VPWR VPWR _08155_ sky130_fd_sc_hd__or2_1
X_10949_ net1816 _05731_ _06165_ VGND VGND VPWR VPWR _06175_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_133_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16456_ _02895_ _03923_ _03924_ _02867_ VGND VGND VPWR VPWR _03925_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13668_ CPU.registerFile\[17\]\[23\] _07404_ VGND VGND VPWR VPWR _08088_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15407_ _08411_ _02892_ _02904_ _07703_ VGND VGND VPWR VPWR _02905_ sky130_fd_sc_hd__a31o_1
X_14590__705 clknet_1_0__leaf__02674_ VGND VGND VPWR VPWR net737 sky130_fd_sc_hd__inv_2
XFILLER_0_26_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12619_ _04654_ _07128_ _07133_ VGND VGND VPWR VPWR _00012_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16387_ CPU.registerFile\[16\]\[28\] _02833_ _02836_ CPU.registerFile\[17\]\[28\]
+ _02764_ VGND VGND VPWR VPWR _03858_ sky130_fd_sc_hd__o221a_1
X_13599_ CPU.registerFile\[13\]\[21\] _07772_ _07773_ CPU.registerFile\[9\]\[21\]
+ _08020_ VGND VGND VPWR VPWR _08021_ sky130_fd_sc_hd__o221a_1
XFILLER_0_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18126_ net189 _02406_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[24\] sky130_fd_sc_hd__dfxtp_1
X_15338_ CPU.registerFile\[18\]\[0\] _02833_ _02836_ CPU.registerFile\[19\]\[0\] _02758_
+ VGND VGND VPWR VPWR _02837_ sky130_fd_sc_hd__o221a_1
XFILLER_0_124_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18057_ net1230 _02337_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_15269_ _02759_ _02762_ _02766_ _02767_ VGND VGND VPWR VPWR _02768_ sky130_fd_sc_hd__a211o_1
X_17008_ net266 _01330_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09830_ _05486_ VGND VGND VPWR VPWR _02510_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410__542 clknet_1_1__leaf__02657_ VGND VGND VPWR VPWR net574 sky130_fd_sc_hd__inv_2
X_09761_ _05449_ VGND VGND VPWR VPWR _02550_ sky130_fd_sc_hd__clkbuf_1
X_08712_ _04325_ _04262_ VGND VGND VPWR VPWR _04432_ sky130_fd_sc_hd__and2b_1
X_09692_ _04758_ _05191_ _04636_ VGND VGND VPWR VPWR _05383_ sky130_fd_sc_hd__mux2_1
Xrebuffer12 net1254 VGND VGND VPWR VPWR net1253 sky130_fd_sc_hd__dlygate4sd1_1
X_08643_ _04230_ _04360_ _04362_ VGND VGND VPWR VPWR _04363_ sky130_fd_sc_hd__o21a_1
Xrebuffer23 net1265 VGND VGND VPWR VPWR net1264 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer34 _04314_ VGND VGND VPWR VPWR net1288 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer45 _04288_ VGND VGND VPWR VPWR net1292 sky130_fd_sc_hd__buf_6
X_14328__469 clknet_1_0__leaf__08465_ VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__inv_2
XFILLER_0_49_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08574_ CPU.instr\[2\] net1275 VGND VGND VPWR VPWR _04294_ sky130_fd_sc_hd__and2b_1
XFILLER_0_89_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09126_ CPU.Jimm\[17\] _04829_ _04831_ VGND VGND VPWR VPWR _04838_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09057_ _04352_ _04210_ _04218_ CPU.aluReg\[25\] VGND VGND VPWR VPWR _04771_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14038__315 clknet_1_0__leaf__08364_ VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__inv_2
Xhold550 CPU.registerFile\[6\]\[7\] VGND VGND VPWR VPWR net1791 sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 CPU.registerFile\[17\]\[19\] VGND VGND VPWR VPWR net1802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 CPU.registerFile\[28\]\[22\] VGND VGND VPWR VPWR net1813 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold583 CPU.registerFile\[12\]\[1\] VGND VGND VPWR VPWR net1824 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold594 CPU.registerFile\[12\]\[23\] VGND VGND VPWR VPWR net1835 sky130_fd_sc_hd__dlygate4sd3_1
X_12769__219 clknet_1_0__leaf__07224_ VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__inv_2
X_14686__791 clknet_1_0__leaf__02684_ VGND VGND VPWR VPWR net823 sky130_fd_sc_hd__inv_2
X_09959_ _05514_ net1624 _05570_ VGND VGND VPWR VPWR _05572_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12970_ _05232_ VGND VGND VPWR VPWR _07411_ sky130_fd_sc_hd__clkbuf_4
Xhold1250 CPU.aluIn1\[30\] VGND VGND VPWR VPWR net2491 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1261 CPU.registerFile\[4\]\[25\] VGND VGND VPWR VPWR net2502 sky130_fd_sc_hd__dlygate4sd3_1
X_11921_ CPU.registerFile\[11\]\[17\] _05700_ _06722_ VGND VGND VPWR VPWR _06727_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1272 CPU.registerFile\[23\]\[14\] VGND VGND VPWR VPWR net2513 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1283 CPU.registerFile\[24\]\[25\] VGND VGND VPWR VPWR net2524 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_401 _02773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1294 CPU.registerFile\[19\]\[18\] VGND VGND VPWR VPWR net2535 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_412 _05070_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14640_ clknet_1_0__leaf__02675_ VGND VGND VPWR VPWR _02680_ sky130_fd_sc_hd__buf_1
X_11852_ _06690_ VGND VGND VPWR VPWR _01642_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_142_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10803_ _06097_ VGND VGND VPWR VPWR _02101_ sky130_fd_sc_hd__clkbuf_1
X_14084__357 clknet_1_1__leaf__08368_ VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__inv_2
X_11783_ net1245 net2124 _06650_ VGND VGND VPWR VPWR _06654_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16310_ CPU.registerFile\[25\]\[26\] CPU.registerFile\[29\]\[26\] _02851_ VGND VGND
+ VPWR VPWR _03783_ sky130_fd_sc_hd__mux2_1
X_13522_ CPU.registerFile\[31\]\[18\] _07629_ _07488_ CPU.registerFile\[27\]\[18\]
+ _07252_ VGND VGND VPWR VPWR _07947_ sky130_fd_sc_hd__o221a_1
XFILLER_0_138_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17290_ net479 _01578_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_527 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10734_ _05541_ net2342 _06056_ VGND VGND VPWR VPWR _06061_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16241_ CPU.registerFile\[7\]\[24\] _03317_ VGND VGND VPWR VPWR _03716_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13453_ CPU.registerFile\[29\]\[16\] _07414_ _07326_ CPU.registerFile\[25\]\[16\]
+ _07489_ VGND VGND VPWR VPWR _07880_ sky130_fd_sc_hd__o221a_1
X_10665_ mapped_spi_flash.state\[3\] _06019_ VGND VGND VPWR VPWR _06022_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_11_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12404_ _07020_ VGND VGND VPWR VPWR _01385_ sky130_fd_sc_hd__clkbuf_1
X_16172_ _03644_ _03648_ _02879_ VGND VGND VPWR VPWR _03649_ sky130_fd_sc_hd__a21o_1
X_13384_ CPU.registerFile\[16\]\[14\] CPU.registerFile\[20\]\[14\] _07648_ VGND VGND
+ VPWR VPWR _07813_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10596_ _05843_ VGND VGND VPWR VPWR _05980_ sky130_fd_sc_hd__buf_2
X_12335_ _04780_ net1786 _06977_ VGND VGND VPWR VPWR _06984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14769__866 clknet_1_0__leaf__02692_ VGND VGND VPWR VPWR net898 sky130_fd_sc_hd__inv_2
X_12266_ CPU.aluReg\[13\] _06934_ _06924_ VGND VGND VPWR VPWR _06935_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_149_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11217_ _06317_ VGND VGND VPWR VPWR _01907_ sky130_fd_sc_hd__clkbuf_1
X_16529__196 clknet_1_1__leaf__03964_ VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__inv_2
X_12197_ net2474 _06881_ _06862_ VGND VGND VPWR VPWR _06882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11148_ CPU.registerFile\[8\]\[5\] _05725_ _06274_ VGND VGND VPWR VPWR _06281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15956_ _03434_ _03438_ _08410_ VGND VGND VPWR VPWR _03439_ sky130_fd_sc_hd__a21o_1
X_11079_ net1696 _05725_ _06237_ VGND VGND VPWR VPWR _06244_ sky130_fd_sc_hd__mux2_1
X_15887_ CPU.registerFile\[9\]\[14\] _02778_ _03125_ VGND VGND VPWR VPWR _03372_ sky130_fd_sc_hd__o21a_1
XFILLER_0_53_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17626_ net815 _01914_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[12\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_82_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17557_ net746 _01845_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17488_ net677 _01776_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16439_ CPU.registerFile\[2\]\[30\] _02872_ _02873_ CPU.registerFile\[3\]\[30\] _05071_
+ VGND VGND VPWR VPWR _03908_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_30_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18109_ net172 _02389_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[7\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_113_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_93_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09813_ net2026 _05253_ _05474_ VGND VGND VPWR VPWR _05478_ sky130_fd_sc_hd__mux2_1
X_16648__92 clknet_1_0__leaf__03989_ VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__inv_2
X_09744_ _04370_ _05431_ _05432_ VGND VGND VPWR VPWR _05433_ sky130_fd_sc_hd__o21a_1
X_09675_ _04418_ _05366_ VGND VGND VPWR VPWR _05367_ sky130_fd_sc_hd__and2b_1
X_15235__144 clknet_1_1__leaf__02754_ VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_38_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08626_ _04245_ _04345_ VGND VGND VPWR VPWR _04346_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_38_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_124_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08557_ _04275_ _04276_ VGND VGND VPWR VPWR _04277_ sky130_fd_sc_hd__or2b_1
XFILLER_0_119_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08488_ CPU.Jimm\[12\] VGND VGND VPWR VPWR _04208_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10450_ _05852_ _04601_ VGND VGND VPWR VPWR _05865_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09109_ CPU.Iimm\[2\] _04496_ _04820_ VGND VGND VPWR VPWR _04821_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10381_ _05812_ _04617_ _04783_ CPU.mem_rstrb VGND VGND VPWR VPWR _05813_ sky130_fd_sc_hd__or4b_2
XFILLER_0_5_690 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12120_ _06832_ VGND VGND VPWR VPWR _01515_ sky130_fd_sc_hd__clkbuf_1
X_12051_ _05008_ net1730 _06794_ VGND VGND VPWR VPWR _06796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold380 CPU.registerFile\[18\]\[29\] VGND VGND VPWR VPWR net1621 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold391 CPU.registerFile\[6\]\[24\] VGND VGND VPWR VPWR net1632 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11002_ _06203_ VGND VGND VPWR VPWR _02008_ sky130_fd_sc_hd__clkbuf_1
X_15810_ _02757_ _03273_ _03283_ _03297_ _02846_ VGND VGND VPWR VPWR _03298_ sky130_fd_sc_hd__a311o_2
XTAP_TAPCELL_ROW_144_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16790_ _04032_ net1568 VGND VGND VPWR VPWR _04101_ sky130_fd_sc_hd__nand2_1
X_15741_ CPU.registerFile\[7\]\[10\] _02806_ _02887_ _03229_ VGND VGND VPWR VPWR _03230_
+ sky130_fd_sc_hd__o211a_1
X_12953_ _04814_ VGND VGND VPWR VPWR _07394_ sky130_fd_sc_hd__clkbuf_4
Xhold1080 CPU.registerFile\[1\]\[16\] VGND VGND VPWR VPWR net2321 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1091 CPU.registerFile\[1\]\[18\] VGND VGND VPWR VPWR net2332 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11904_ net2174 _05683_ _06711_ VGND VGND VPWR VPWR _06718_ sky130_fd_sc_hd__mux2_1
X_15672_ CPU.registerFile\[15\]\[8\] CPU.registerFile\[11\]\[8\] _02773_ VGND VGND
+ VPWR VPWR _03163_ sky130_fd_sc_hd__mux2_1
X_12884_ _07237_ VGND VGND VPWR VPWR _07326_ sky130_fd_sc_hd__clkbuf_8
XANTENNA_220 clknet_1_0__leaf__02749_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_231 clknet_1_1__leaf__07219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13949__235 clknet_1_0__leaf__07226_ VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__inv_2
XANTENNA_242 _03064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17411_ net600 _01699_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[4\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_253 _05045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11835_ _06681_ VGND VGND VPWR VPWR _01650_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_264 _05129_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_275 _05543_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_25_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_286 _05710_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17342_ net531 _01630_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[6\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_297 _07271_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11766_ _04762_ net1756 _06639_ VGND VGND VPWR VPWR _06645_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ _07392_ _07925_ _07929_ _07232_ VGND VGND VPWR VPWR _07930_ sky130_fd_sc_hd__o211a_2
X_17273_ net462 _01561_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_60_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10717_ _05524_ net2129 _06045_ VGND VGND VPWR VPWR _06052_ sky130_fd_sc_hd__mux2_1
X_14485_ clknet_1_1__leaf__02664_ VGND VGND VPWR VPWR _02665_ sky130_fd_sc_hd__buf_1
XFILLER_0_71_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11697_ mapped_spi_ram.rcv_data\[12\] _06601_ VGND VGND VPWR VPWR _06602_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16224_ CPU.registerFile\[12\]\[24\] _03118_ VGND VGND VPWR VPWR _03699_ sky130_fd_sc_hd__or2_1
X_13436_ net1533 _07229_ _07863_ _07135_ VGND VGND VPWR VPWR _01310_ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10648_ mapped_spi_flash.rcv_data\[0\] _05969_ VGND VGND VPWR VPWR _06009_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer3 _04547_ VGND VGND VPWR VPWR net1285 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_130_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16155_ CPU.aluIn1\[21\] _03081_ _03631_ _03632_ VGND VGND VPWR VPWR _02435_ sky130_fd_sc_hd__o211a_1
X_16590__61 clknet_1_1__leaf__03970_ VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__inv_2
XFILLER_0_12_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_13367_ _07296_ _07796_ VGND VGND VPWR VPWR _07797_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10579_ mapped_spi_flash.rcv_data\[31\] _05970_ VGND VGND VPWR VPWR _05971_ sky130_fd_sc_hd__or2_1
X_14357__495 clknet_1_0__leaf__08468_ VGND VGND VPWR VPWR net527 sky130_fd_sc_hd__inv_2
X_15106_ net1465 _07191_ VGND VGND VPWR VPWR _02740_ sky130_fd_sc_hd__nand2_1
X_12318_ _04412_ _06856_ _06973_ VGND VGND VPWR VPWR _06974_ sky130_fd_sc_hd__a21oi_1
X_16086_ CPU.registerFile\[5\]\[20\] CPU.registerFile\[4\]\[20\] _05092_ VGND VGND
+ VPWR VPWR _03565_ sky130_fd_sc_hd__mux2_1
X_13298_ CPU.registerFile\[15\]\[11\] _07629_ _07488_ CPU.registerFile\[11\]\[11\]
+ _07252_ VGND VGND VPWR VPWR _07730_ sky130_fd_sc_hd__o221a_1
X_13995__277 clknet_1_0__leaf__08359_ VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__inv_2
X_12249_ _06921_ VGND VGND VPWR VPWR _01441_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_75_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16988_ clknet_leaf_28_clk _01314_ VGND VGND VPWR VPWR CPU.rs2\[19\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_147_Right_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_917 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15939_ CPU.registerFile\[22\]\[15\] _03032_ VGND VGND VPWR VPWR _03423_ sky130_fd_sc_hd__and2_1
X_09460_ _04434_ _05160_ VGND VGND VPWR VPWR _05161_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_35_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14067__341 clknet_1_1__leaf__08367_ VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_35_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14522__643 clknet_1_1__leaf__02668_ VGND VGND VPWR VPWR net675 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_106_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17609_ net798 _01897_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[27\] sky130_fd_sc_hd__dfxtp_1
X_09391_ _04845_ _04897_ VGND VGND VPWR VPWR _05095_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_16_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_59_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_688 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_116_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_839 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_126_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_114_Right_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14605__718 clknet_1_0__leaf__02676_ VGND VGND VPWR VPWR net750 sky130_fd_sc_hd__inv_2
X_09727_ CPU.aluIn1\[0\] _04302_ VGND VGND VPWR VPWR _05417_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_2_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09658_ _04420_ _05350_ VGND VGND VPWR VPWR _05351_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14798__892 clknet_1_0__leaf__02695_ VGND VGND VPWR VPWR net924 sky130_fd_sc_hd__inv_2
X_08609_ CPU.aluIn1\[14\] _04257_ VGND VGND VPWR VPWR _04329_ sky130_fd_sc_hd__nand2_1
X_09589_ _05283_ VGND VGND VPWR VPWR _05284_ sky130_fd_sc_hd__buf_6
XFILLER_0_139_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14497__620 clknet_1_0__leaf__02666_ VGND VGND VPWR VPWR net652 sky130_fd_sc_hd__inv_2
X_11620_ mapped_spi_ram.snd_bitcount\[3\] _06549_ VGND VGND VPWR VPWR _06550_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11551_ net1409 _06495_ _06503_ _06006_ VGND VGND VPWR VPWR _01755_ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10502_ _04516_ _04542_ _04515_ VGND VGND VPWR VPWR _05909_ sky130_fd_sc_hd__a21oi_1
X_14270_ _04683_ _04740_ _05433_ VGND VGND VPWR VPWR _08449_ sky130_fd_sc_hd__mux2_1
X_11482_ _06458_ VGND VGND VPWR VPWR _01783_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_502 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13221_ CPU.registerFile\[21\]\[9\] _07403_ _07619_ CPU.registerFile\[17\]\[9\] _07250_
+ VGND VGND VPWR VPWR _07655_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_21_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10433_ _05852_ _04588_ VGND VGND VPWR VPWR _05853_ sky130_fd_sc_hd__nor2_1
X_13152_ CPU.registerFile\[29\]\[7\] _07325_ _07326_ CPU.registerFile\[25\]\[7\] _07249_
+ VGND VGND VPWR VPWR _07588_ sky130_fd_sc_hd__o221a_1
X_10364_ _05541_ net2341 _05799_ VGND VGND VPWR VPWR _05804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12103_ _06823_ VGND VGND VPWR VPWR _01523_ sky130_fd_sc_hd__clkbuf_1
X_13083_ _07238_ VGND VGND VPWR VPWR _07521_ sky130_fd_sc_hd__buf_4
X_17960_ net1148 _02244_ VGND VGND VPWR VPWR CPU.registerFile\[21\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_10295_ _05541_ net2322 _05762_ VGND VGND VPWR VPWR _05767_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12034_ _04731_ net2127 _06783_ VGND VGND VPWR VPWR _06787_ sky130_fd_sc_hd__mux2_1
X_16911_ CPU.mem_wdata\[1\] _04180_ _04184_ _04176_ VGND VGND VPWR VPWR _02639_ sky130_fd_sc_hd__o211a_1
X_17891_ net1080 _02175_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[9\] sky130_fd_sc_hd__dfxtp_1
X_16842_ _03977_ _04138_ VGND VGND VPWR VPWR _04139_ sky130_fd_sc_hd__nand2b_4
XTAP_TAPCELL_ROW_70_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16627__73 clknet_1_1__leaf__03971_ VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__inv_2
X_16773_ _04027_ _04039_ _05022_ VGND VGND VPWR VPWR _04087_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12936_ CPU.registerFile\[3\]\[2\] _07373_ _07375_ _07376_ VGND VGND VPWR VPWR _07377_
+ sky130_fd_sc_hd__o211a_1
X_15724_ _03015_ _03211_ _03213_ _03019_ VGND VGND VPWR VPWR _03214_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16642__87 clknet_1_0__leaf__03988_ VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__inv_2
X_15655_ CPU.registerFile\[5\]\[7\] CPU.registerFile\[4\]\[7\] _03146_ VGND VGND VPWR
+ VPWR _03147_ sky130_fd_sc_hd__mux2_1
X_12867_ _07230_ _07270_ _07307_ _07309_ VGND VGND VPWR VPWR _07310_ sky130_fd_sc_hd__a211o_1
X_11818_ _05426_ net2137 _06638_ VGND VGND VPWR VPWR _06672_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_157_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15586_ _06515_ VGND VGND VPWR VPWR _03080_ sky130_fd_sc_hd__buf_2
XFILLER_0_157_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12798_ CPU.registerFile\[18\]\[0\] CPU.registerFile\[22\]\[0\] _07240_ VGND VGND
+ VPWR VPWR _07241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17325_ net514 _01613_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11749_ mapped_spi_ram.rcv_bitcount\[0\] net13 VGND VGND VPWR VPWR _06635_ sky130_fd_sc_hd__and2b_1
Xclkbuf_1_1__f__03963_ clknet_0__03963_ VGND VGND VPWR VPWR clknet_1_1__leaf__03963_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_44_839 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17256_ net446 _01544_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13419_ _07844_ _07846_ _04972_ VGND VGND VPWR VPWR _07847_ sky130_fd_sc_hd__mux2_1
X_16207_ _03681_ _03682_ _02875_ VGND VGND VPWR VPWR _03683_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_77_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17187_ clknet_leaf_29_clk _01475_ VGND VGND VPWR VPWR CPU.Jimm\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16138_ _03611_ _03615_ _03138_ VGND VGND VPWR VPWR _03616_ sky130_fd_sc_hd__a21o_1
XFILLER_0_141_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08960_ _04678_ VGND VGND VPWR VPWR _04679_ sky130_fd_sc_hd__clkbuf_4
X_16069_ _03195_ _03546_ _03547_ _03548_ _03245_ VGND VGND VPWR VPWR _03549_ sky130_fd_sc_hd__a221o_1
XFILLER_0_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_5_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_90_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08891_ CPU.PC\[18\] _04586_ _04609_ _04610_ VGND VGND VPWR VPWR _04611_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_108_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09512_ _05210_ VGND VGND VPWR VPWR _02560_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_88_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09443_ _04436_ _05144_ VGND VGND VPWR VPWR _05145_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_121_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_09374_ _04333_ _04392_ _04440_ VGND VGND VPWR VPWR _05079_ sky130_fd_sc_hd__or3_1
XFILLER_0_148_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13978__261 clknet_1_1__leaf__08358_ VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__inv_2
XFILLER_0_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10080_ net2185 _04731_ _05633_ VGND VGND VPWR VPWR _05637_ sky130_fd_sc_hd__mux2_1
X_13770_ _07653_ _08185_ _08186_ VGND VGND VPWR VPWR _08187_ sky130_fd_sc_hd__o21ai_1
X_10982_ net1586 _05696_ _06190_ VGND VGND VPWR VPWR _06193_ sky130_fd_sc_hd__mux2_1
X_12721_ _07179_ _07202_ VGND VGND VPWR VPWR _07203_ sky130_fd_sc_hd__nor2_4
XFILLER_0_78_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15440_ CPU.registerFile\[7\]\[2\] _05092_ VGND VGND VPWR VPWR _02937_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_26_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12652_ CPU.cycles\[13\] CPU.cycles\[14\] _07150_ VGND VGND VPWR VPWR _07152_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_26_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_139_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11603_ net1350 _06524_ _06540_ _06539_ VGND VGND VPWR VPWR _01740_ sky130_fd_sc_hd__o211a_1
X_15371_ CPU.registerFile\[1\]\[1\] _02867_ _02868_ _08405_ VGND VGND VPWR VPWR _02869_
+ sky130_fd_sc_hd__a22o_1
X_12583_ net1995 _05358_ _07107_ VGND VGND VPWR VPWR _07115_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17110_ clknet_leaf_14_clk _00043_ VGND VGND VPWR VPWR CPU.cycles\[6\] sky130_fd_sc_hd__dfxtp_1
X_18090_ net153 _02370_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_11534_ _05816_ net1321 _06489_ _06492_ net1313 VGND VGND VPWR VPWR _01761_ sky130_fd_sc_hd__a32o_1
XFILLER_0_20_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_885 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17041_ net299 _01363_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_152_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11465_ _06449_ VGND VGND VPWR VPWR _01791_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13204_ _05284_ VGND VGND VPWR VPWR _07638_ sky130_fd_sc_hd__buf_4
X_10416_ _05840_ VGND VGND VPWR VPWR _02230_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11396_ _05520_ net2218 _06408_ VGND VGND VPWR VPWR _06413_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__02661_ _02661_ VGND VGND VPWR VPWR clknet_0__02661_ sky130_fd_sc_hd__clkbuf_16
X_13135_ CPU.registerFile\[18\]\[7\] CPU.registerFile\[22\]\[7\] _07233_ VGND VGND
+ VPWR VPWR _07571_ sky130_fd_sc_hd__mux2_1
X_10347_ _05524_ net1810 _05788_ VGND VGND VPWR VPWR _05795_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17943_ net1132 _02227_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[23\] sky130_fd_sc_hd__dfxtp_1
X_13066_ CPU.registerFile\[21\]\[5\] _07502_ _07503_ CPU.registerFile\[17\]\[5\] _07300_
+ VGND VGND VPWR VPWR _07504_ sky130_fd_sc_hd__o221a_1
X_10278_ _05524_ net2210 _05751_ VGND VGND VPWR VPWR _05758_ sky130_fd_sc_hd__mux2_1
X_12017_ _06777_ VGND VGND VPWR VPWR _01564_ sky130_fd_sc_hd__clkbuf_1
X_17874_ net1063 _02158_ VGND VGND VPWR VPWR mapped_spi_flash.clk_div sky130_fd_sc_hd__dfxtp_1
X_14469__596 clknet_1_1__leaf__02662_ VGND VGND VPWR VPWR net628 sky130_fd_sc_hd__inv_2
X_16825_ _04115_ _04126_ per_uart.uart0.tx_bitcount\[0\] VGND VGND VPWR VPWR _04127_
+ sky130_fd_sc_hd__mux2_1
X_16756_ _04052_ _05087_ _04006_ VGND VGND VPWR VPWR _04073_ sky130_fd_sc_hd__or3b_1
XFILLER_0_88_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15707_ CPU.registerFile\[11\]\[9\] _02861_ VGND VGND VPWR VPWR _03197_ sky130_fd_sc_hd__or2_1
XFILLER_0_158_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12919_ _07359_ VGND VGND VPWR VPWR _07360_ sky130_fd_sc_hd__buf_4
X_13899_ _07818_ _08310_ _08311_ VGND VGND VPWR VPWR _08312_ sky130_fd_sc_hd__o21a_1
X_16687_ _04589_ VGND VGND VPWR VPWR _04015_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_103_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15638_ _05406_ VGND VGND VPWR VPWR _03130_ sky130_fd_sc_hd__buf_4
XPHY_EDGE_ROW_14_Left_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18357_ clknet_leaf_4_clk _02635_ VGND VGND VPWR VPWR per_uart.uart0.rx_ack sky130_fd_sc_hd__dfxtp_1
X_15569_ _03059_ _03060_ _03062_ _02945_ VGND VGND VPWR VPWR _03063_ sky130_fd_sc_hd__o22a_1
XFILLER_0_56_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17308_ net497 _01596_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_09090_ _04462_ _04801_ VGND VGND VPWR VPWR _04802_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18288_ net121 _02568_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_142_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14634__744 clknet_1_1__leaf__02679_ VGND VGND VPWR VPWR net776 sky130_fd_sc_hd__inv_2
XFILLER_0_153_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17239_ net429 _01527_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold902 CPU.registerFile\[28\]\[9\] VGND VGND VPWR VPWR net2143 sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 CPU.registerFile\[1\]\[21\] VGND VGND VPWR VPWR net2154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold924 CPU.registerFile\[19\]\[5\] VGND VGND VPWR VPWR net2165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold935 CPU.registerFile\[2\]\[11\] VGND VGND VPWR VPWR net2176 sky130_fd_sc_hd__dlygate4sd3_1
Xhold946 CPU.registerFile\[13\]\[7\] VGND VGND VPWR VPWR net2187 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold957 CPU.registerFile\[14\]\[14\] VGND VGND VPWR VPWR net2198 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__08435_ _08435_ VGND VGND VPWR VPWR clknet_0__08435_ sky130_fd_sc_hd__clkbuf_16
Xhold968 CPU.registerFile\[3\]\[10\] VGND VGND VPWR VPWR net2209 sky130_fd_sc_hd__dlygate4sd3_1
X_09992_ _05547_ net2223 _05581_ VGND VGND VPWR VPWR _05589_ sky130_fd_sc_hd__mux2_1
Xhold979 CPU.registerFile\[31\]\[17\] VGND VGND VPWR VPWR net2220 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_23_Left_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__08366_ _08366_ VGND VGND VPWR VPWR clknet_0__08366_ sky130_fd_sc_hd__clkbuf_16
X_08943_ CPU.Bimm\[3\] VGND VGND VPWR VPWR _04663_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_4_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08874_ _04506_ _04582_ _04588_ _04593_ VGND VGND VPWR VPWR _04594_ sky130_fd_sc_hd__o211ai_4
X_14959__1037 clknet_1_1__leaf__02711_ VGND VGND VPWR VPWR net1069 sky130_fd_sc_hd__inv_2
X_14680__786 clknet_1_0__leaf__02683_ VGND VGND VPWR VPWR net818 sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_32_Left_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09426_ _05114_ _05115_ _05123_ _05128_ VGND VGND VPWR VPWR _05129_ sky130_fd_sc_hd__or4b_4
XFILLER_0_137_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14717__819 clknet_1_1__leaf__02687_ VGND VGND VPWR VPWR net851 sky130_fd_sc_hd__inv_2
X_09357_ _04841_ _04901_ VGND VGND VPWR VPWR _05063_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09288_ _04960_ _04996_ VGND VGND VPWR VPWR _04997_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11250_ _06323_ VGND VGND VPWR VPWR _06335_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_132_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10201_ _05169_ VGND VGND VPWR VPWR _05710_ sky130_fd_sc_hd__clkbuf_4
X_11181_ _06298_ VGND VGND VPWR VPWR _01924_ sky130_fd_sc_hd__clkbuf_1
X_10132_ net1945 _05381_ _05655_ VGND VGND VPWR VPWR _05664_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14940_ clknet_1_0__leaf__02708_ VGND VGND VPWR VPWR _02710_ sky130_fd_sc_hd__buf_1
X_10063_ net1983 _05381_ _05618_ VGND VGND VPWR VPWR _05627_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__03966_ clknet_0__03966_ VGND VGND VPWR VPWR clknet_1_0__leaf__03966_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_50_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16610_ _03980_ VGND VGND VPWR VPWR _02542_ sky130_fd_sc_hd__clkbuf_1
X_13822_ CPU.registerFile\[13\]\[28\] _07772_ _07773_ CPU.registerFile\[9\]\[28\]
+ _08236_ VGND VGND VPWR VPWR _08237_ sky130_fd_sc_hd__o221a_1
X_17590_ net779 _01878_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13753_ CPU.registerFile\[15\]\[25\] CPU.registerFile\[7\]\[25\] _04648_ VGND VGND
+ VPWR VPWR _08171_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10965_ net1607 _05679_ _06179_ VGND VGND VPWR VPWR _06184_ sky130_fd_sc_hd__mux2_1
X_12704_ net1466 _07185_ VGND VGND VPWR VPWR _07186_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13684_ CPU.registerFile\[14\]\[23\] CPU.registerFile\[10\]\[23\] _07399_ VGND VGND
+ VPWR VPWR _08104_ sky130_fd_sc_hd__mux2_1
X_16472_ _03227_ _03938_ _03939_ _03030_ VGND VGND VPWR VPWR _03940_ sky130_fd_sc_hd__a22o_1
X_10896_ _06147_ VGND VGND VPWR VPWR _02058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18211_ net52 _02491_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_12635_ net1462 _07140_ VGND VGND VPWR VPWR _07143_ sky130_fd_sc_hd__nor2_1
X_15423_ CPU.registerFile\[28\]\[2\] _05049_ VGND VGND VPWR VPWR _02920_ sky130_fd_sc_hd__or2_1
XFILLER_0_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_122_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18142_ clknet_leaf_19_clk _02422_ VGND VGND VPWR VPWR CPU.aluIn1\[8\] sky130_fd_sc_hd__dfxtp_2
X_15354_ _02851_ VGND VGND VPWR VPWR _02852_ sky130_fd_sc_hd__clkbuf_8
X_12566_ net2412 _05169_ _07096_ VGND VGND VPWR VPWR _07106_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11517_ _06480_ VGND VGND VPWR VPWR _01766_ sky130_fd_sc_hd__clkbuf_1
X_15285_ _05361_ VGND VGND VPWR VPWR _02784_ sky130_fd_sc_hd__clkbuf_4
X_18073_ net136 _02353_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_12497_ _07069_ VGND VGND VPWR VPWR _01341_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17024_ net282 _01346_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[18\] sky130_fd_sc_hd__dfxtp_1
X_14236_ clknet_1_1__leaf__08433_ VGND VGND VPWR VPWR _08434_ sky130_fd_sc_hd__buf_1
Xhold209 mapped_spi_ram.rcv_data\[30\] VGND VGND VPWR VPWR net1450 sky130_fd_sc_hd__dlygate4sd3_1
X_11448_ _06440_ VGND VGND VPWR VPWR _01799_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__02713_ _02713_ VGND VGND VPWR VPWR clknet_0__02713_ sky130_fd_sc_hd__clkbuf_16
X_14167_ _08420_ VGND VGND VPWR VPWR _01484_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11379_ _05503_ net2524 _06397_ VGND VGND VPWR VPWR _06404_ sky130_fd_sc_hd__mux2_1
X_13118_ _07554_ VGND VGND VPWR VPWR _07555_ sky130_fd_sc_hd__buf_4
X_14098_ _08372_ _08374_ _08376_ VGND VGND VPWR VPWR _08377_ sky130_fd_sc_hd__and3_1
X_13049_ _07237_ VGND VGND VPWR VPWR _07488_ sky130_fd_sc_hd__buf_4
X_17926_ net1115 _02210_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14215__391 clknet_1_1__leaf__08431_ VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__inv_2
X_17857_ net1046 _02141_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_16808_ net2 _07200_ VGND VGND VPWR VPWR _04115_ sky130_fd_sc_hd__and2_1
X_16498__168 clknet_1_0__leaf__02756_ VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__inv_2
X_08590_ _04285_ _04287_ _04307_ _04309_ VGND VGND VPWR VPWR _04310_ sky130_fd_sc_hd__a31o_1
X_17788_ net977 _02072_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_85_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16739_ _03995_ _05143_ _07132_ VGND VGND VPWR VPWR _04059_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09211_ CPU.PC\[13\] CPU.PC\[12\] _04922_ VGND VGND VPWR VPWR _04923_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09142_ CPU.PC\[11\] _04853_ VGND VGND VPWR VPWR _04854_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09073_ _04782_ _04785_ net1277 VGND VGND VPWR VPWR _04786_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold710 CPU.registerFile\[2\]\[23\] VGND VGND VPWR VPWR net1951 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_685 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold721 CPU.registerFile\[31\]\[31\] VGND VGND VPWR VPWR net1962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 CPU.registerFile\[31\]\[12\] VGND VGND VPWR VPWR net1973 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold743 CPU.registerFile\[15\]\[30\] VGND VGND VPWR VPWR net1984 sky130_fd_sc_hd__dlygate4sd3_1
Xhold754 CPU.registerFile\[4\]\[4\] VGND VGND VPWR VPWR net1995 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold765 CPU.registerFile\[24\]\[29\] VGND VGND VPWR VPWR net2006 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold776 CPU.registerFile\[31\]\[10\] VGND VGND VPWR VPWR net2017 sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 CPU.registerFile\[21\]\[14\] VGND VGND VPWR VPWR net2028 sky130_fd_sc_hd__dlygate4sd3_1
X_09975_ _05530_ net1646 _05570_ VGND VGND VPWR VPWR _05580_ sky130_fd_sc_hd__mux2_1
Xhold798 CPU.registerFile\[15\]\[17\] VGND VGND VPWR VPWR net2039 sky130_fd_sc_hd__dlygate4sd3_1
X_08926_ mapped_spi_ram.rcv_data\[31\] net17 _04618_ mapped_spi_flash.rcv_data\[31\]
+ VGND VGND VPWR VPWR _04646_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08857_ CPU.aluIn1\[21\] _04495_ VGND VGND VPWR VPWR _04577_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_28_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__02702_ clknet_0__02702_ VGND VGND VPWR VPWR clknet_1_0__leaf__02702_
+ sky130_fd_sc_hd__clkbuf_16
X_08788_ CPU.aluIn1\[12\] CPU.Bimm\[12\] VGND VGND VPWR VPWR _04508_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10750_ _05557_ _06032_ VGND VGND VPWR VPWR _06069_ sky130_fd_sc_hd__nand2_2
XFILLER_0_138_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14305__448 clknet_1_0__leaf__08463_ VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__inv_2
X_09409_ _04215_ _04621_ VGND VGND VPWR VPWR _05112_ sky130_fd_sc_hd__nand2_2
X_10681_ _04665_ _04663_ _04664_ CPU.writeBack VGND VGND VPWR VPWR _06032_ sky130_fd_sc_hd__and4_2
XFILLER_0_48_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12420_ net1244 net2220 _07024_ VGND VGND VPWR VPWR _07029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12351_ _06992_ VGND VGND VPWR VPWR _01410_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11302_ _05495_ net2164 _06360_ VGND VGND VPWR VPWR _06363_ sky130_fd_sc_hd__mux2_1
X_12282_ CPU.aluIn1\[9\] _06946_ _06927_ VGND VGND VPWR VPWR _06947_ sky130_fd_sc_hd__mux2_1
X_11233_ _06326_ VGND VGND VPWR VPWR _01900_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_52_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11164_ _05493_ net2334 _06288_ VGND VGND VPWR VPWR _06290_ sky130_fd_sc_hd__mux2_1
X_10115_ _05632_ VGND VGND VPWR VPWR _05655_ sky130_fd_sc_hd__buf_4
X_11095_ _06253_ VGND VGND VPWR VPWR _01965_ sky130_fd_sc_hd__clkbuf_1
X_15972_ CPU.registerFile\[20\]\[16\] CPU.registerFile\[21\]\[16\] _08394_ VGND VGND
+ VPWR VPWR _03455_ sky130_fd_sc_hd__mux2_1
X_17711_ net900 _00009_ VGND VGND VPWR VPWR mapped_spi_ram.state\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_147_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10046_ _05595_ VGND VGND VPWR VPWR _05618_ sky130_fd_sc_hd__buf_4
X_14663__770 clknet_1_0__leaf__02682_ VGND VGND VPWR VPWR net802 sky130_fd_sc_hd__inv_2
Xhold70 _06621_ VGND VGND VPWR VPWR net1311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 mapped_spi_ram.rcv_data\[25\] VGND VGND VPWR VPWR net1322 sky130_fd_sc_hd__dlygate4sd3_1
X_17642_ net831 _01930_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[28\] sky130_fd_sc_hd__dfxtp_1
Xhold92 _00008_ VGND VGND VPWR VPWR net1333 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13805_ CPU.registerFile\[15\]\[27\] _07236_ _07239_ CPU.registerFile\[11\]\[27\]
+ _07820_ VGND VGND VPWR VPWR _08221_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_67_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17573_ net762 _01861_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11997_ _05150_ net1619 _06758_ VGND VGND VPWR VPWR _06767_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10948_ _06174_ VGND VGND VPWR VPWR _02033_ sky130_fd_sc_hd__clkbuf_1
X_13736_ CPU.registerFile\[13\]\[25\] CPU.registerFile\[12\]\[25\] _04985_ VGND VGND
+ VPWR VPWR _08154_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16455_ CPU.registerFile\[19\]\[30\] CPU.registerFile\[17\]\[30\] _03025_ VGND VGND
+ VPWR VPWR _03924_ sky130_fd_sc_hd__mux2_1
X_10879_ _06137_ VGND VGND VPWR VPWR _02065_ sky130_fd_sc_hd__clkbuf_1
X_13667_ _08081_ _08083_ _08085_ _08086_ VGND VGND VPWR VPWR _08087_ sky130_fd_sc_hd__o22a_1
XFILLER_0_144_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14061__336 clknet_1_1__leaf__08366_ VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_80_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15406_ _02867_ _02893_ _02902_ _02903_ VGND VGND VPWR VPWR _02904_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_14_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12618_ CPU.state\[3\] _07133_ VGND VGND VPWR VPWR _00014_ sky130_fd_sc_hd__nor2_1
X_13598_ _07260_ _08019_ VGND VGND VPWR VPWR _08020_ sky130_fd_sc_hd__or2_1
X_16386_ CPU.registerFile\[20\]\[28\] CPU.registerFile\[21\]\[28\] _08395_ VGND VGND
+ VPWR VPWR _03857_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18125_ net188 _02405_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[23\] sky130_fd_sc_hd__dfxtp_1
X_12549_ _07097_ VGND VGND VPWR VPWR _01284_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14958__1036 clknet_1_1__leaf__02711_ VGND VGND VPWR VPWR net1068 sky130_fd_sc_hd__inv_2
X_15337_ _02835_ VGND VGND VPWR VPWR _02836_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_112_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18056_ net1229 _02336_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[18\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_1 CPU.Bimm\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15268_ _08396_ VGND VGND VPWR VPWR _02767_ sky130_fd_sc_hd__buf_4
X_17007_ net265 _01329_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14746__845 clknet_1_1__leaf__02690_ VGND VGND VPWR VPWR net877 sky130_fd_sc_hd__inv_2
X_09760_ net1770 _05448_ _04667_ VGND VGND VPWR VPWR _05449_ sky130_fd_sc_hd__mux2_1
X_08711_ _04399_ _04320_ VGND VGND VPWR VPWR _04431_ sky130_fd_sc_hd__nand2_1
X_16506__175 clknet_1_1__leaf__03962_ VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__inv_2
X_17909_ net1098 net1469 VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[27\] sky130_fd_sc_hd__dfxtp_1
X_09691_ _05382_ VGND VGND VPWR VPWR _02553_ sky130_fd_sc_hd__clkbuf_1
X_08642_ _04228_ _04361_ VGND VGND VPWR VPWR _04362_ sky130_fd_sc_hd__nor2_1
Xrebuffer13 net1255 VGND VGND VPWR VPWR net1254 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer24 net1266 VGND VGND VPWR VPWR net1265 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_96_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer35 _04517_ VGND VGND VPWR VPWR net1276 sky130_fd_sc_hd__dlymetal6s4s_1
Xrebuffer46 _04415_ VGND VGND VPWR VPWR net1293 sky130_fd_sc_hd__dlygate4sd1_1
X_08573_ CPU.instr\[3\] _04291_ _04292_ VGND VGND VPWR VPWR _04293_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_77_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14792__887 clknet_1_1__leaf__02694_ VGND VGND VPWR VPWR net919 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_33_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09125_ CPU.PC\[18\] _04836_ VGND VGND VPWR VPWR _04837_ sky130_fd_sc_hd__and2_1
X_14491__615 clknet_1_0__leaf__02665_ VGND VGND VPWR VPWR net647 sky130_fd_sc_hd__inv_2
XFILLER_0_127_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_98_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09056_ _04234_ _04683_ VGND VGND VPWR VPWR _04770_ sky130_fd_sc_hd__nor2_1
Xhold540 CPU.registerFile\[30\]\[1\] VGND VGND VPWR VPWR net1781 sky130_fd_sc_hd__dlygate4sd3_1
Xhold551 CPU.registerFile\[13\]\[25\] VGND VGND VPWR VPWR net1792 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_694 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold562 CPU.registerFile\[19\]\[28\] VGND VGND VPWR VPWR net1803 sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 CPU.registerFile\[4\]\[20\] VGND VGND VPWR VPWR net1814 sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 per_uart.uart0.rxd_reg\[7\] VGND VGND VPWR VPWR net1825 sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 CPU.registerFile\[27\]\[15\] VGND VGND VPWR VPWR net1836 sky130_fd_sc_hd__dlygate4sd3_1
X_14231__406 clknet_1_0__leaf__08432_ VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__inv_2
X_09958_ _05571_ VGND VGND VPWR VPWR _02467_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_129_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08909_ _04506_ VGND VGND VPWR VPWR _04629_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_129_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09889_ _05527_ VGND VGND VPWR VPWR _02492_ sky130_fd_sc_hd__clkbuf_1
Xhold1240 CPU.PC\[21\] VGND VGND VPWR VPWR net2481 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1251 CPU.registerFile\[1\]\[12\] VGND VGND VPWR VPWR net2492 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1262 CPU.aluReg\[17\] VGND VGND VPWR VPWR net2503 sky130_fd_sc_hd__dlygate4sd3_1
X_11920_ _06726_ VGND VGND VPWR VPWR _01610_ sky130_fd_sc_hd__clkbuf_1
Xhold1273 CPU.aluReg\[26\] VGND VGND VPWR VPWR net2514 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1284 CPU.registerFile\[16\]\[14\] VGND VGND VPWR VPWR net2525 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1295 CPU.registerFile\[11\]\[21\] VGND VGND VPWR VPWR net2536 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_402 _02773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11851_ net2167 _05698_ _06686_ VGND VGND VPWR VPWR _06690_ sky130_fd_sc_hd__mux2_1
XANTENNA_413 _05333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10802_ _05541_ net2303 _06092_ VGND VGND VPWR VPWR _06097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11782_ _06653_ VGND VGND VPWR VPWR _01675_ sky130_fd_sc_hd__clkbuf_1
X_15212__123 clknet_1_0__leaf__02752_ VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__inv_2
XFILLER_0_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13521_ CPU.registerFile\[30\]\[18\] CPU.registerFile\[26\]\[18\] _07399_ VGND VGND
+ VPWR VPWR _07946_ sky130_fd_sc_hd__mux2_1
X_10733_ _06060_ VGND VGND VPWR VPWR _02134_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13452_ CPU.registerFile\[28\]\[16\] CPU.registerFile\[24\]\[16\] _07476_ VGND VGND
+ VPWR VPWR _07879_ sky130_fd_sc_hd__mux2_1
X_16240_ _03710_ _03714_ _03138_ VGND VGND VPWR VPWR _03715_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_62_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10664_ _05850_ _06019_ _06021_ net1320 VGND VGND VPWR VPWR _02164_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_11_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12403_ _04780_ net2097 _07013_ VGND VGND VPWR VPWR _07020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16171_ _02924_ _03645_ _03646_ _03647_ _02930_ VGND VGND VPWR VPWR _03648_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13383_ CPU.registerFile\[23\]\[14\] _07282_ _07811_ VGND VGND VPWR VPWR _07812_
+ sky130_fd_sc_hd__o21ai_2
X_10595_ mapped_spi_flash.rcv_data\[23\] _05970_ VGND VGND VPWR VPWR _05979_ sky130_fd_sc_hd__or2_1
X_12334_ _06983_ VGND VGND VPWR VPWR _01418_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15053_ clknet_1_1__leaf__02720_ VGND VGND VPWR VPWR _02722_ sky130_fd_sc_hd__buf_1
X_12265_ CPU.aluIn1\[13\] _06933_ _06927_ VGND VGND VPWR VPWR _06934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_128_Right_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11216_ _05545_ net2237 _06310_ VGND VGND VPWR VPWR _06317_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12196_ CPU.aluIn1\[29\] _06880_ _06865_ VGND VGND VPWR VPWR _06881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11147_ _06280_ VGND VGND VPWR VPWR _01940_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15955_ _02771_ _03435_ _03436_ _03437_ _02807_ VGND VGND VPWR VPWR _03438_ sky130_fd_sc_hd__a221o_1
X_11078_ _06243_ VGND VGND VPWR VPWR _01972_ sky130_fd_sc_hd__clkbuf_1
X_14906_ clknet_1_1__leaf__02697_ VGND VGND VPWR VPWR _02706_ sky130_fd_sc_hd__buf_1
X_10029_ _05609_ VGND VGND VPWR VPWR _02402_ sky130_fd_sc_hd__clkbuf_1
X_15886_ CPU.registerFile\[13\]\[14\] _03123_ VGND VGND VPWR VPWR _03371_ sky130_fd_sc_hd__or2_1
X_17625_ net814 _01913_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[11\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_19_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17556_ net745 _01844_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13719_ _07330_ _08137_ VGND VGND VPWR VPWR _08138_ sky130_fd_sc_hd__or2_1
X_15187__100 clknet_1_1__leaf__02750_ VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__inv_2
X_17487_ net676 _01775_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_16438_ CPU.registerFile\[6\]\[30\] CPU.registerFile\[7\]\[30\] _02870_ VGND VGND
+ VPWR VPWR _03907_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16369_ CPU.registerFile\[28\]\[28\] _03064_ VGND VGND VPWR VPWR _03840_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18108_ net171 _02388_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18039_ net1212 _02319_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14334__474 clknet_1_1__leaf__08466_ VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__inv_2
XFILLER_0_10_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09812_ _05477_ VGND VGND VPWR VPWR _02519_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13972__256 clknet_1_0__leaf__08357_ VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__inv_2
X_09743_ _04369_ _04207_ VGND VGND VPWR VPWR _05432_ sky130_fd_sc_hd__or2_1
X_09674_ _04417_ _04408_ _04416_ VGND VGND VPWR VPWR _05366_ sky130_fd_sc_hd__or3_1
X_08625_ CPU.aluIn1\[20\] _04246_ _04344_ VGND VGND VPWR VPWR _04345_ sky130_fd_sc_hd__a21o_1
XFILLER_0_96_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_6_Left_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_124_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08556_ CPU.aluIn1\[6\] _04274_ VGND VGND VPWR VPWR _04276_ sky130_fd_sc_hd__or2_1
X_14800__894 clknet_1_1__leaf__02695_ VGND VGND VPWR VPWR net926 sky130_fd_sc_hd__inv_2
XFILLER_0_65_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08487_ CPU.rs2\[31\] _04201_ _04206_ VGND VGND VPWR VPWR _04207_ sky130_fd_sc_hd__a21o_1
XFILLER_0_147_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14044__320 clknet_1_0__leaf__08365_ VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__inv_2
XFILLER_0_92_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12775__224 clknet_1_1__leaf__07225_ VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__inv_2
XFILLER_0_123_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09108_ _04819_ VGND VGND VPWR VPWR _04820_ sky130_fd_sc_hd__buf_2
XFILLER_0_122_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10380_ net1418 VGND VGND VPWR VPWR _05812_ sky130_fd_sc_hd__inv_2
X_14417__549 clknet_1_0__leaf__02657_ VGND VGND VPWR VPWR net581 sky130_fd_sc_hd__inv_2
X_09039_ _04671_ _04751_ _04753_ _04678_ VGND VGND VPWR VPWR _04754_ sky130_fd_sc_hd__o211a_1
X_12050_ _06795_ VGND VGND VPWR VPWR _01548_ sky130_fd_sc_hd__clkbuf_1
Xhold370 CPU.registerFile\[6\]\[30\] VGND VGND VPWR VPWR net1611 sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 CPU.registerFile\[2\]\[0\] VGND VGND VPWR VPWR net1622 sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ net2298 _05715_ _06201_ VGND VGND VPWR VPWR _06203_ sky130_fd_sc_hd__mux2_1
Xhold392 CPU.registerFile\[30\]\[12\] VGND VGND VPWR VPWR net1633 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_144_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15740_ CPU.registerFile\[6\]\[10\] _02819_ VGND VGND VPWR VPWR _03229_ sky130_fd_sc_hd__or2_1
X_12952_ _07360_ _07386_ _07391_ _07392_ VGND VGND VPWR VPWR _07393_ sky130_fd_sc_hd__o211a_1
X_14957__1035 clknet_1_1__leaf__02711_ VGND VGND VPWR VPWR net1067 sky130_fd_sc_hd__inv_2
Xhold1070 CPU.registerFile\[6\]\[5\] VGND VGND VPWR VPWR net2311 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 CPU.registerFile\[20\]\[7\] VGND VGND VPWR VPWR net2322 sky130_fd_sc_hd__dlygate4sd3_1
X_11903_ _06717_ VGND VGND VPWR VPWR _01618_ sky130_fd_sc_hd__clkbuf_1
Xhold1092 CPU.registerFile\[19\]\[16\] VGND VGND VPWR VPWR net2333 sky130_fd_sc_hd__dlygate4sd3_1
X_15671_ _02759_ _03159_ _03161_ _02767_ VGND VGND VPWR VPWR _03162_ sky130_fd_sc_hd__a211o_1
X_15179__1204 clknet_1_0__leaf__02748_ VGND VGND VPWR VPWR net1236 sky130_fd_sc_hd__inv_2
XANTENNA_210 _07914_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12883_ _07234_ VGND VGND VPWR VPWR _07325_ sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_47_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_221 clknet_1_1__leaf__02750_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_305 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_232 CPU.mem_wdata\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17410_ net599 _01698_ VGND VGND VPWR VPWR mapped_spi_ram.rcv_data\[3\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_243 _03064_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_254 _05045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11834_ net1644 _05681_ _06675_ VGND VGND VPWR VPWR _06681_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_265 _05333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_276 _05551_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17341_ net530 _01629_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[5\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_287 _05719_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_298 _07318_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11765_ _06644_ VGND VGND VPWR VPWR _01683_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14775__871 clknet_1_0__leaf__02693_ VGND VGND VPWR VPWR net903 sky130_fd_sc_hd__inv_2
XFILLER_0_67_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ _06051_ VGND VGND VPWR VPWR _02142_ sky130_fd_sc_hd__clkbuf_1
X_13504_ _07288_ _07928_ VGND VGND VPWR VPWR _07929_ sky130_fd_sc_hd__or2_1
X_17272_ net461 _01560_ VGND VGND VPWR VPWR CPU.registerFile\[12\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_14484_ clknet_1_1__leaf__07222_ VGND VGND VPWR VPWR _02664_ sky130_fd_sc_hd__buf_1
X_11696_ _06576_ VGND VGND VPWR VPWR _06601_ sky130_fd_sc_hd__clkbuf_2
X_16223_ CPU.registerFile\[14\]\[24\] CPU.registerFile\[10\]\[24\] _02787_ VGND VGND
+ VPWR VPWR _03698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_114_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13435_ _07230_ _07848_ _07862_ _07309_ VGND VGND VPWR VPWR _07863_ sky130_fd_sc_hd__a211o_1
X_10647_ net2268 _05967_ _06008_ _06006_ VGND VGND VPWR VPWR _02167_ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer4 net1287 VGND VGND VPWR VPWR net1286 sky130_fd_sc_hd__clkbuf_2
X_13366_ CPU.registerFile\[30\]\[13\] CPU.registerFile\[26\]\[13\] _04938_ VGND VGND
+ VPWR VPWR _07796_ sky130_fd_sc_hd__mux2_1
X_16154_ _06515_ VGND VGND VPWR VPWR _03632_ sky130_fd_sc_hd__buf_4
X_10578_ _05969_ VGND VGND VPWR VPWR _05970_ sky130_fd_sc_hd__buf_2
XFILLER_0_134_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15105_ _07191_ _02739_ _02727_ VGND VGND VPWR VPWR _02282_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12317_ CPU.aluReg\[1\] _06872_ _06856_ VGND VGND VPWR VPWR _06973_ sky130_fd_sc_hd__a21oi_1
X_13297_ CPU.registerFile\[14\]\[11\] CPU.registerFile\[10\]\[11\] _07399_ VGND VGND
+ VPWR VPWR _07729_ sky130_fd_sc_hd__mux2_1
X_16085_ CPU.aluIn1\[19\] _02958_ _03545_ _03564_ _02995_ VGND VGND VPWR VPWR _02433_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_121_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12248_ net2503 _06920_ _06891_ VGND VGND VPWR VPWR _06921_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12179_ CPU.aluShamt\[1\] CPU.aluShamt\[0\] VGND VGND VPWR VPWR _06868_ sky130_fd_sc_hd__and2_1
X_16987_ clknet_leaf_28_clk _01313_ VGND VGND VPWR VPWR CPU.rs2\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15938_ CPU.registerFile\[21\]\[15\] CPU.registerFile\[23\]\[15\] _02769_ VGND VGND
+ VPWR VPWR _03422_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_15869_ CPU.registerFile\[1\]\[13\] _02939_ _03354_ _02943_ VGND VGND VPWR VPWR _03355_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_35_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14858__946 clknet_1_1__leaf__02701_ VGND VGND VPWR VPWR net978 sky130_fd_sc_hd__inv_2
X_17608_ net797 _01896_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[26\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_35_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09390_ _04782_ _05093_ _04622_ _04681_ VGND VGND VPWR VPWR _05094_ sky130_fd_sc_hd__a22oi_2
XTAP_TAPCELL_ROW_106_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17539_ net728 _01827_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_745 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_126_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09726_ _05415_ _04413_ VGND VGND VPWR VPWR _05416_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09657_ _04419_ _04407_ _04418_ VGND VGND VPWR VPWR _05350_ sky130_fd_sc_hd__nor3_1
XFILLER_0_97_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08608_ _04326_ _04260_ _04327_ VGND VGND VPWR VPWR _04328_ sky130_fd_sc_hd__a21o_1
X_09588_ _05282_ VGND VGND VPWR VPWR _05283_ sky130_fd_sc_hd__buf_8
XFILLER_0_96_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08539_ CPU.rs2\[13\] _04199_ _04204_ VGND VGND VPWR VPWR _04259_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11550_ net1394 _06499_ _06489_ _06502_ VGND VGND VPWR VPWR _06503_ sky130_fd_sc_hd__a211o_1
XFILLER_0_37_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10501_ net1366 _05892_ _05908_ _05885_ VGND VGND VPWR VPWR _02213_ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11481_ _05537_ net2449 _06455_ VGND VGND VPWR VPWR _06458_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13220_ CPU.registerFile\[16\]\[9\] CPU.registerFile\[20\]\[9\] _07258_ VGND VGND
+ VPWR VPWR _07654_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10432_ _05817_ VGND VGND VPWR VPWR _05852_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_137_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13151_ CPU.registerFile\[28\]\[7\] CPU.registerFile\[24\]\[7\] _07476_ VGND VGND
+ VPWR VPWR _07587_ sky130_fd_sc_hd__mux2_1
X_10363_ _05803_ VGND VGND VPWR VPWR _02247_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12102_ _04731_ net2058 _06819_ VGND VGND VPWR VPWR _06823_ sky130_fd_sc_hd__mux2_1
X_13082_ CPU.registerFile\[8\]\[5\] CPU.registerFile\[12\]\[5\] _07318_ VGND VGND
+ VPWR VPWR _07520_ sky130_fd_sc_hd__mux2_1
X_10294_ _05766_ VGND VGND VPWR VPWR _02294_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_57_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12033_ _06786_ VGND VGND VPWR VPWR _01556_ sky130_fd_sc_hd__clkbuf_1
X_16910_ net1637 _04182_ VGND VGND VPWR VPWR _04184_ sky130_fd_sc_hd__or2_1
X_13955__240 clknet_1_0__leaf__08356_ VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__inv_2
X_17890_ net1079 _02174_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16841_ per_uart.uart0.uart_rxd2 _04137_ _03975_ VGND VGND VPWR VPWR _04138_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_69_Left_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14016__296 clknet_1_0__leaf__08361_ VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__inv_2
X_16772_ _04032_ net1691 VGND VGND VPWR VPWR _04086_ sky130_fd_sc_hd__nand2_1
X_15723_ _02796_ _03212_ VGND VGND VPWR VPWR _03213_ sky130_fd_sc_hd__or2_1
X_12935_ _04938_ VGND VGND VPWR VPWR _07376_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_125_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15654_ net15 VGND VGND VPWR VPWR _03146_ sky130_fd_sc_hd__buf_4
XFILLER_0_157_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12866_ _07308_ VGND VGND VPWR VPWR _07309_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_68_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11817_ _06671_ VGND VGND VPWR VPWR _01658_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18373_ net41 net32 VGND VGND VPWR VPWR mapped_spi_ram.div_counter\[5\] sky130_fd_sc_hd__dfxtp_1
X_15585_ _02757_ _03045_ _03056_ _03078_ _02846_ VGND VGND VPWR VPWR _03079_ sky130_fd_sc_hd__a311o_1
XFILLER_0_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12797_ _05282_ VGND VGND VPWR VPWR _07240_ sky130_fd_sc_hd__buf_4
XFILLER_0_56_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17324_ net513 _01612_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_1__f__03962_ clknet_0__03962_ VGND VGND VPWR VPWR clknet_1_1__leaf__03962_
+ sky130_fd_sc_hd__clkbuf_16
X_11748_ net1349 _06627_ net13 _06634_ VGND VGND VPWR VPWR _01690_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Left_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17255_ net445 _01543_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_11679_ net1478 _06588_ VGND VGND VPWR VPWR _06592_ sky130_fd_sc_hd__or2_1
XFILLER_0_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16206_ CPU.registerFile\[8\]\[23\] CPU.registerFile\[12\]\[23\] _02798_ VGND VGND
+ VPWR VPWR _03682_ sky130_fd_sc_hd__mux2_1
X_13418_ CPU.registerFile\[1\]\[15\] _07255_ _07845_ _07318_ VGND VGND VPWR VPWR _07846_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17186_ clknet_leaf_29_clk _01474_ VGND VGND VPWR VPWR CPU.Jimm\[16\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_77_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_737 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16137_ _02885_ _03612_ _03613_ _03614_ _03022_ VGND VGND VPWR VPWR _03615_ sky130_fd_sc_hd__a221o_1
X_13349_ CPU.registerFile\[2\]\[13\] CPU.registerFile\[3\]\[13\] _07263_ VGND VGND
+ VPWR VPWR _07779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_901 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16068_ CPU.registerFile\[10\]\[19\] _02816_ _02910_ VGND VGND VPWR VPWR _03548_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_90_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_781 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08890_ _04590_ _04605_ VGND VGND VPWR VPWR _04610_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_87_Left_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09511_ net1737 _05209_ _05189_ VGND VGND VPWR VPWR _05210_ sky130_fd_sc_hd__mux2_1
X_14446__575 clknet_1_0__leaf__02660_ VGND VGND VPWR VPWR net607 sky130_fd_sc_hd__inv_2
X_09442_ _04435_ _04398_ _04434_ VGND VGND VPWR VPWR _05144_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_88_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14184__363 clknet_1_1__leaf__08428_ VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_121_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09373_ _04334_ _05077_ VGND VGND VPWR VPWR _05078_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_96_Left_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_615 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_144_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14912__995 clknet_1_0__leaf__02706_ VGND VGND VPWR VPWR net1027 sky130_fd_sc_hd__inv_2
X_14956__1034 clknet_1_0__leaf__02711_ VGND VGND VPWR VPWR net1066 sky130_fd_sc_hd__inv_2
XFILLER_0_43_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15178__1203 clknet_1_1__leaf__02748_ VGND VGND VPWR VPWR net1235 sky130_fd_sc_hd__inv_2
X_14611__723 clknet_1_0__leaf__02677_ VGND VGND VPWR VPWR net755 sky130_fd_sc_hd__inv_2
XFILLER_0_112_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09709_ CPU.PC\[2\] _04955_ _05390_ _04974_ _05399_ VGND VGND VPWR VPWR _05400_ sky130_fd_sc_hd__o221ai_2
X_10981_ _06192_ VGND VGND VPWR VPWR _02018_ sky130_fd_sc_hd__clkbuf_1
X_12720_ _07200_ _07201_ VGND VGND VPWR VPWR _07202_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12651_ net1514 _07150_ VGND VGND VPWR VPWR _00019_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_26_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_155_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11602_ net1392 _06517_ _06496_ CPU.mem_wdata\[7\] _06508_ VGND VGND VPWR VPWR _06540_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_139_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15370_ CPU.registerFile\[5\]\[1\] CPU.registerFile\[4\]\[1\] _02806_ VGND VGND VPWR
+ VPWR _02868_ sky130_fd_sc_hd__mux2_1
X_12582_ _07114_ VGND VGND VPWR VPWR _01268_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11533_ _05816_ net1327 _06489_ _06492_ net1321 VGND VGND VPWR VPWR _01762_ sky130_fd_sc_hd__a32o_1
XFILLER_0_136_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17040_ net298 _01362_ VGND VGND VPWR VPWR CPU.registerFile\[31\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_11464_ _05520_ net1996 _06444_ VGND VGND VPWR VPWR _06449_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_152_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13203_ CPU.registerFile\[5\]\[9\] CPU.registerFile\[4\]\[9\] _07262_ VGND VGND VPWR
+ VPWR _07637_ sky130_fd_sc_hd__mux2_1
X_10415_ _05830_ _05839_ VGND VGND VPWR VPWR _05840_ sky130_fd_sc_hd__and2_1
XFILLER_0_151_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_11395_ _06412_ VGND VGND VPWR VPWR _01824_ sky130_fd_sc_hd__clkbuf_1
X_14887__972 clknet_1_1__leaf__02704_ VGND VGND VPWR VPWR net1004 sky130_fd_sc_hd__inv_2
XFILLER_0_150_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13134_ _07300_ VGND VGND VPWR VPWR _07570_ sky130_fd_sc_hd__buf_4
Xclkbuf_0__02660_ _02660_ VGND VGND VPWR VPWR clknet_0__02660_ sky130_fd_sc_hd__clkbuf_16
X_10346_ _05794_ VGND VGND VPWR VPWR _02255_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_72_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13065_ _07238_ VGND VGND VPWR VPWR _07503_ sky130_fd_sc_hd__buf_4
X_17942_ net1131 _02226_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[22\] sky130_fd_sc_hd__dfxtp_1
X_10277_ _05757_ VGND VGND VPWR VPWR _02302_ sky130_fd_sc_hd__clkbuf_1
X_12016_ _05359_ net2263 _06769_ VGND VGND VPWR VPWR _06777_ sky130_fd_sc_hd__mux2_1
X_17873_ net1062 _02157_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16824_ _07178_ net20 _04192_ VGND VGND VPWR VPWR _04126_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16755_ _04027_ _04039_ _05085_ VGND VGND VPWR VPWR _04072_ sky130_fd_sc_hd__a21o_1
X_15706_ CPU.registerFile\[9\]\[9\] CPU.registerFile\[13\]\[9\] _02999_ VGND VGND
+ VPWR VPWR _03196_ sky130_fd_sc_hd__mux2_1
X_12918_ _04785_ VGND VGND VPWR VPWR _07359_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16686_ _08457_ _04011_ _04012_ _04013_ VGND VGND VPWR VPWR _04014_ sky130_fd_sc_hd__a31o_1
XFILLER_0_158_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13898_ CPU.registerFile\[15\]\[30\] _07236_ _07239_ CPU.registerFile\[11\]\[30\]
+ _07820_ VGND VGND VPWR VPWR _08311_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_103_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15637_ CPU.registerFile\[30\]\[7\] CPU.registerFile\[26\]\[7\] _02787_ VGND VGND
+ VPWR VPWR _03129_ sky130_fd_sc_hd__mux2_1
X_12849_ _04935_ VGND VGND VPWR VPWR _07292_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_158_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18356_ clknet_leaf_1_clk net1312 VGND VGND VPWR VPWR per_uart.uart0.uart_rxd2 sky130_fd_sc_hd__dfxtp_1
X_15568_ CPU.registerFile\[1\]\[5\] _02814_ _03061_ _02943_ VGND VGND VPWR VPWR _03062_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17307_ net496 _01595_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18287_ net120 _02567_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15499_ _05843_ VGND VGND VPWR VPWR _02995_ sky130_fd_sc_hd__buf_2
XFILLER_0_127_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_823 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17238_ net428 _01526_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold903 CPU.registerFile\[10\]\[28\] VGND VGND VPWR VPWR net2144 sky130_fd_sc_hd__dlygate4sd3_1
X_17169_ clknet_leaf_25_clk _01457_ VGND VGND VPWR VPWR CPU.mem_wmask\[1\] sky130_fd_sc_hd__dfxtp_1
Xhold914 CPU.registerFile\[20\]\[31\] VGND VGND VPWR VPWR net2155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold925 CPU.registerFile\[25\]\[24\] VGND VGND VPWR VPWR net2166 sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 CPU.registerFile\[24\]\[5\] VGND VGND VPWR VPWR net2177 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__08434_ _08434_ VGND VGND VPWR VPWR clknet_0__08434_ sky130_fd_sc_hd__clkbuf_16
Xhold947 CPU.registerFile\[20\]\[11\] VGND VGND VPWR VPWR net2188 sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 CPU.registerFile\[23\]\[28\] VGND VGND VPWR VPWR net2199 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09991_ _05588_ VGND VGND VPWR VPWR _02451_ sky130_fd_sc_hd__clkbuf_1
Xhold969 CPU.registerFile\[20\]\[15\] VGND VGND VPWR VPWR net2210 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__08365_ _08365_ VGND VGND VPWR VPWR clknet_0__08365_ sky130_fd_sc_hd__clkbuf_16
X_08942_ _04660_ _04661_ VGND VGND VPWR VPWR _04662_ sky130_fd_sc_hd__or2_4
Xclkbuf_1_1__f__02689_ clknet_0__02689_ VGND VGND VPWR VPWR clknet_1_1__leaf__02689_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_4_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08873_ CPU.PC\[23\] _04586_ _04592_ VGND VGND VPWR VPWR _04593_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09425_ _04818_ _05125_ _05127_ _04916_ VGND VGND VPWR VPWR _05128_ sky130_fd_sc_hd__o22a_1
XFILLER_0_94_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09356_ CPU.PC\[17\] _04925_ VGND VGND VPWR VPWR _05062_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_09287_ _04343_ _04385_ _04449_ VGND VGND VPWR VPWR _04996_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10200_ _05709_ VGND VGND VPWR VPWR _02331_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11180_ _05509_ net1968 _06288_ VGND VGND VPWR VPWR _06298_ sky130_fd_sc_hd__mux2_1
X_10131_ _05663_ VGND VGND VPWR VPWR _02354_ sky130_fd_sc_hd__clkbuf_1
X_10062_ _05626_ VGND VGND VPWR VPWR _02386_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__03965_ clknet_0__03965_ VGND VGND VPWR VPWR clknet_1_0__leaf__03965_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_50_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13821_ _07370_ _08235_ VGND VGND VPWR VPWR _08236_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_832 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13752_ CPU.registerFile\[11\]\[25\] CPU.registerFile\[3\]\[25\] _04648_ VGND VGND
+ VPWR VPWR _08170_ sky130_fd_sc_hd__mux2_1
X_10964_ _06183_ VGND VGND VPWR VPWR _02026_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12703_ per_uart.uart0.enable16_counter\[6\] _07184_ VGND VGND VPWR VPWR _07185_
+ sky130_fd_sc_hd__or2_1
X_16471_ CPU.registerFile\[19\]\[31\] CPU.registerFile\[17\]\[31\] _02874_ VGND VGND
+ VPWR VPWR _03939_ sky130_fd_sc_hd__mux2_1
X_13683_ _08099_ _08102_ _07305_ VGND VGND VPWR VPWR _08103_ sky130_fd_sc_hd__a21o_1
X_10895_ net1570 _05677_ _06143_ VGND VGND VPWR VPWR _06147_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18210_ net51 _02490_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_442 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15422_ CPU.registerFile\[30\]\[2\] CPU.registerFile\[26\]\[2\] _02918_ VGND VGND
+ VPWR VPWR _02919_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_902 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12634_ CPU.cycles\[6\] _07140_ VGND VGND VPWR VPWR _07142_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18141_ clknet_leaf_19_clk _02421_ VGND VGND VPWR VPWR CPU.aluIn1\[7\] sky130_fd_sc_hd__dfxtp_2
XFILLER_0_93_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15353_ _05405_ VGND VGND VPWR VPWR _02851_ sky130_fd_sc_hd__clkbuf_8
X_12565_ _07105_ VGND VGND VPWR VPWR _01276_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18072_ net135 _02352_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_11516_ _05830_ net2529 _06031_ VGND VGND VPWR VPWR _06480_ sky130_fd_sc_hd__and3_1
X_15284_ _02771_ _02774_ _02776_ _02781_ _02782_ VGND VGND VPWR VPWR _02783_ sky130_fd_sc_hd__a221o_1
X_12496_ net1942 _05708_ _07060_ VGND VGND VPWR VPWR _07069_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17023_ net281 _01345_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_14235_ clknet_1_0__leaf__07222_ VGND VGND VPWR VPWR _08433_ sky130_fd_sc_hd__buf_1
XFILLER_0_150_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11447_ _05503_ net2113 _06433_ VGND VGND VPWR VPWR _06440_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__02712_ _02712_ VGND VGND VPWR VPWR clknet_0__02712_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11378_ _06403_ VGND VGND VPWR VPWR _01832_ sky130_fd_sc_hd__clkbuf_1
X_14166_ CPU.Bimm\[6\] _04758_ _08413_ VGND VGND VPWR VPWR _08420_ sky130_fd_sc_hd__mux2_1
X_13117_ _04971_ VGND VGND VPWR VPWR _07554_ sky130_fd_sc_hd__buf_4
X_10329_ _05785_ VGND VGND VPWR VPWR _02263_ sky130_fd_sc_hd__clkbuf_1
X_14097_ _04716_ net1273 VGND VGND VPWR VPWR _08376_ sky130_fd_sc_hd__nand2_1
X_13048_ CPU.registerFile\[8\]\[4\] CPU.registerFile\[12\]\[4\] _07265_ VGND VGND
+ VPWR VPWR _07487_ sky130_fd_sc_hd__mux2_1
X_17925_ net1114 _02209_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_147_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17856_ net1045 _02140_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[14\] sky130_fd_sc_hd__dfxtp_1
X_16807_ net2222 per_uart.tx_busy VGND VGND VPWR VPWR _04114_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17787_ net976 _02071_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14955__1033 clknet_1_0__leaf__02711_ VGND VGND VPWR VPWR net1065 sky130_fd_sc_hd__inv_2
X_16738_ _04052_ _05138_ _04006_ VGND VGND VPWR VPWR _04058_ sky130_fd_sc_hd__or3b_1
XFILLER_0_72_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15177__1202 clknet_1_0__leaf__02748_ VGND VGND VPWR VPWR net1234 sky130_fd_sc_hd__inv_2
X_16669_ _08436_ _08459_ _05377_ VGND VGND VPWR VPWR _03999_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09210_ CPU.PC\[11\] _04921_ VGND VGND VPWR VPWR _04922_ sky130_fd_sc_hd__and2_1
XFILLER_0_146_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_902 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09141_ _04499_ CPU.Iimm\[0\] _04661_ _04830_ VGND VGND VPWR VPWR _04853_ sky130_fd_sc_hd__a22o_1
X_18339_ clknet_leaf_4_clk _02619_ VGND VGND VPWR VPWR per_uart.rx_data\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14558__676 clknet_1_0__leaf__02671_ VGND VGND VPWR VPWR net708 sky130_fd_sc_hd__inv_2
XFILLER_0_72_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09072_ mapped_spi_ram.rcv_data\[0\] _04783_ _04784_ mapped_spi_flash.rcv_data\[0\]
+ VGND VGND VPWR VPWR _04785_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_112_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold700 CPU.registerFile\[20\]\[27\] VGND VGND VPWR VPWR net1941 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold711 CPU.registerFile\[22\]\[17\] VGND VGND VPWR VPWR net1952 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold722 CPU.registerFile\[17\]\[1\] VGND VGND VPWR VPWR net1963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold733 per_uart.d_in_uart\[3\] VGND VGND VPWR VPWR net1974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 CPU.registerFile\[1\]\[3\] VGND VGND VPWR VPWR net1985 sky130_fd_sc_hd__dlygate4sd3_1
Xhold755 CPU.registerFile\[25\]\[17\] VGND VGND VPWR VPWR net1996 sky130_fd_sc_hd__dlygate4sd3_1
Xhold766 CPU.registerFile\[18\]\[31\] VGND VGND VPWR VPWR net2007 sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 CPU.registerFile\[12\]\[28\] VGND VGND VPWR VPWR net2018 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 CPU.registerFile\[26\]\[1\] VGND VGND VPWR VPWR net2029 sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ _05579_ VGND VGND VPWR VPWR _02459_ sky130_fd_sc_hd__clkbuf_1
Xhold799 CPU.registerFile\[26\]\[22\] VGND VGND VPWR VPWR net2040 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_08925_ _04594_ _04599_ _04613_ VGND VGND VPWR VPWR _04645_ sky130_fd_sc_hd__nor3_2
X_08856_ CPU.aluIn1\[21\] _04495_ VGND VGND VPWR VPWR _04576_ sky130_fd_sc_hd__nor2_1
X_14723__824 clknet_1_0__leaf__02688_ VGND VGND VPWR VPWR net856 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__02701_ clknet_0__02701_ VGND VGND VPWR VPWR clknet_1_0__leaf__02701_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08787_ CPU.aluIn1\[12\] CPU.Bimm\[12\] VGND VGND VPWR VPWR _04507_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09408_ mapped_spi_ram.rcv_data\[22\] _04689_ _04691_ mapped_spi_flash.rcv_data\[22\]
+ VGND VGND VPWR VPWR _05111_ sky130_fd_sc_hd__a22o_1
X_10680_ _06030_ net1315 VGND VGND VPWR VPWR _02158_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09339_ _05045_ VGND VGND VPWR VPWR _05046_ sky130_fd_sc_hd__buf_12
XFILLER_0_62_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_109_Right_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_117_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12350_ net1245 net1848 _06988_ VGND VGND VPWR VPWR _06992_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11301_ _06362_ VGND VGND VPWR VPWR _01868_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12281_ CPU.aluReg\[10\] CPU.aluReg\[8\] _06939_ VGND VGND VPWR VPWR _06946_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11232_ net1760 _05673_ _06324_ VGND VGND VPWR VPWR _06326_ sky130_fd_sc_hd__mux2_1
X_14020_ clknet_1_0__leaf__07223_ VGND VGND VPWR VPWR _08362_ sky130_fd_sc_hd__buf_1
XFILLER_0_120_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11163_ _06289_ VGND VGND VPWR VPWR _01933_ sky130_fd_sc_hd__clkbuf_1
X_10114_ _05654_ VGND VGND VPWR VPWR _02362_ sky130_fd_sc_hd__clkbuf_1
X_15971_ _03450_ _03451_ _03453_ _02945_ VGND VGND VPWR VPWR _03454_ sky130_fd_sc_hd__o22a_2
X_11094_ net1557 _05668_ _06252_ VGND VGND VPWR VPWR _06253_ sky130_fd_sc_hd__mux2_1
X_17710_ net899 net1333 VGND VGND VPWR VPWR mapped_spi_ram.state\[0\] sky130_fd_sc_hd__dfxtp_1
X_10045_ _05617_ VGND VGND VPWR VPWR _02394_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold71 per_uart.uart0.uart_rxd1 VGND VGND VPWR VPWR net1312 sky130_fd_sc_hd__dlygate4sd3_1
X_17641_ net830 _01929_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[27\] sky130_fd_sc_hd__dfxtp_1
Xhold82 _01721_ VGND VGND VPWR VPWR net1323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 mapped_spi_ram.snd_bitcount\[3\] VGND VGND VPWR VPWR net1334 sky130_fd_sc_hd__dlygate4sd3_1
X_13804_ CPU.registerFile\[14\]\[27\] CPU.registerFile\[10\]\[27\] _07480_ VGND VGND
+ VPWR VPWR _08220_ sky130_fd_sc_hd__mux2_1
X_17572_ net761 _01860_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_14784_ clknet_1_1__leaf__02686_ VGND VGND VPWR VPWR _02694_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_67_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11996_ _06766_ VGND VGND VPWR VPWR _01574_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_67_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13735_ CPU.registerFile\[8\]\[25\] CPU.registerFile\[9\]\[25\] _05338_ VGND VGND
+ VPWR VPWR _08153_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10947_ net1584 _05729_ _06165_ VGND VGND VPWR VPWR _06174_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_100_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16597__68 clknet_1_0__leaf__03970_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__inv_2
XFILLER_0_42_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16454_ _03921_ _03922_ _02898_ VGND VGND VPWR VPWR _03923_ sky130_fd_sc_hd__mux2_1
X_13666_ CPU.registerFile\[29\]\[23\] _08082_ _07256_ CPU.registerFile\[25\]\[23\]
+ _07405_ VGND VGND VPWR VPWR _08086_ sky130_fd_sc_hd__a221o_1
X_10878_ net1681 _05729_ _06128_ VGND VGND VPWR VPWR _06137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15405_ _05384_ VGND VGND VPWR VPWR _02903_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_14_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12617_ _07132_ _04589_ CPU.state\[2\] CPU.state\[0\] VGND VGND VPWR VPWR _07133_
+ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_14_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16385_ _02827_ _03854_ _03855_ VGND VGND VPWR VPWR _03856_ sky130_fd_sc_hd__o21ai_1
X_13597_ CPU.registerFile\[8\]\[21\] CPU.registerFile\[12\]\[21\] _07233_ VGND VGND
+ VPWR VPWR _08019_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__07219_ clknet_0__07219_ VGND VGND VPWR VPWR clknet_1_0__leaf__07219_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_143_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18124_ net187 _02404_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[22\] sky130_fd_sc_hd__dfxtp_1
X_15336_ _02834_ VGND VGND VPWR VPWR _02835_ sky130_fd_sc_hd__buf_4
X_12548_ net1895 _04981_ _07096_ VGND VGND VPWR VPWR _07097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18055_ net1228 _02335_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[17\] sky130_fd_sc_hd__dfxtp_1
X_15267_ CPU.registerFile\[8\]\[0\] _02763_ _02764_ _02765_ VGND VGND VPWR VPWR _02766_
+ sky130_fd_sc_hd__o211a_1
X_12479_ _07048_ VGND VGND VPWR VPWR _07060_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_2 CPU.Iimm\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17006_ net264 _01328_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14149_ _05361_ VGND VGND VPWR VPWR _08410_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_158_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08710_ _04429_ _04402_ _04266_ VGND VGND VPWR VPWR _04430_ sky130_fd_sc_hd__o21a_1
X_17908_ net1097 net1405 VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[26\] sky130_fd_sc_hd__dfxtp_1
X_09690_ net1817 _05381_ _05189_ VGND VGND VPWR VPWR _05382_ sky130_fd_sc_hd__mux2_1
X_08641_ CPU.aluIn1\[28\] _04227_ VGND VGND VPWR VPWR _04361_ sky130_fd_sc_hd__nor2_1
X_17839_ net1028 _02123_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[29\] sky130_fd_sc_hd__dfxtp_1
Xrebuffer14 net1256 VGND VGND VPWR VPWR net1255 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer25 net1267 VGND VGND VPWR VPWR net1266 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer36 _04543_ VGND VGND VPWR VPWR net1289 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer47 _04415_ VGND VGND VPWR VPWR net1294 sky130_fd_sc_hd__dlygate4sd1_1
X_08572_ CPU.instr\[4\] VGND VGND VPWR VPWR _04292_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_507 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_119_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15159__1186 clknet_1_1__leaf__02746_ VGND VGND VPWR VPWR net1218 sky130_fd_sc_hd__inv_2
XFILLER_0_8_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_754 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_288 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09124_ CPU.Jimm\[18\] _04829_ _04831_ VGND VGND VPWR VPWR _04836_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09055_ _04672_ _04765_ _04767_ _04768_ VGND VGND VPWR VPWR _04769_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_131_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold530 CPU.registerFile\[24\]\[20\] VGND VGND VPWR VPWR net1771 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold541 CPU.registerFile\[12\]\[25\] VGND VGND VPWR VPWR net1782 sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 CPU.registerFile\[5\]\[4\] VGND VGND VPWR VPWR net1793 sky130_fd_sc_hd__dlygate4sd3_1
Xhold563 CPU.registerFile\[30\]\[9\] VGND VGND VPWR VPWR net1804 sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 CPU.registerFile\[25\]\[1\] VGND VGND VPWR VPWR net1815 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold585 CPU.registerFile\[26\]\[15\] VGND VGND VPWR VPWR net1826 sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 CPU.registerFile\[13\]\[13\] VGND VGND VPWR VPWR net1837 sky130_fd_sc_hd__dlygate4sd3_1
X_09957_ _05511_ net1718 _05570_ VGND VGND VPWR VPWR _05571_ sky130_fd_sc_hd__mux2_1
X_14311__453 clknet_1_0__leaf__08464_ VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__inv_2
X_08908_ _04522_ _04533_ _04627_ VGND VGND VPWR VPWR _04628_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_129_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ _05526_ net1998 _05512_ VGND VGND VPWR VPWR _05527_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_129_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1230 mapped_spi_ram.rcv_data\[9\] VGND VGND VPWR VPWR net2471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1241 CPU.registerFile\[24\]\[24\] VGND VGND VPWR VPWR net2482 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1252 CPU.registerFile\[23\]\[5\] VGND VGND VPWR VPWR net2493 sky130_fd_sc_hd__dlygate4sd3_1
X_08839_ CPU.aluIn1\[16\] _04494_ VGND VGND VPWR VPWR _04559_ sky130_fd_sc_hd__nand2_1
Xhold1263 mapped_spi_ram.rcv_bitcount\[1\] VGND VGND VPWR VPWR net2504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1274 CPU.registerFile\[15\]\[5\] VGND VGND VPWR VPWR net2515 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1285 CPU.registerFile\[22\]\[25\] VGND VGND VPWR VPWR net2526 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1296 CPU.registerFile\[11\]\[4\] VGND VGND VPWR VPWR net2537 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_403 _03138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11850_ _06689_ VGND VGND VPWR VPWR _01643_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_414 _05333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_142_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ _06096_ VGND VGND VPWR VPWR _02102_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11781_ _05027_ net2080 _06650_ VGND VGND VPWR VPWR _06653_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13520_ _07411_ _07941_ _07944_ VGND VGND VPWR VPWR _07945_ sky130_fd_sc_hd__or3_1
XFILLER_0_83_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10732_ _05539_ net2315 _06056_ VGND VGND VPWR VPWR _06060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13451_ _07870_ _07877_ _07395_ VGND VGND VPWR VPWR _07878_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_62_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10663_ _06018_ _06020_ VGND VGND VPWR VPWR _06021_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12402_ _07019_ VGND VGND VPWR VPWR _01386_ sky130_fd_sc_hd__clkbuf_1
X_16170_ CPU.registerFile\[25\]\[22\] _02943_ _02860_ VGND VGND VPWR VPWR _03647_
+ sky130_fd_sc_hd__o21a_1
X_10594_ net1704 _05968_ _05978_ _05936_ VGND VGND VPWR VPWR _02190_ sky130_fd_sc_hd__o211a_1
X_13382_ CPU.registerFile\[19\]\[14\] _07618_ _07810_ _07417_ _07253_ VGND VGND VPWR
+ VPWR _07811_ sky130_fd_sc_hd__o221a_1
XFILLER_0_63_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12333_ _04762_ net1902 _06977_ VGND VGND VPWR VPWR _06983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12264_ CPU.aluReg\[14\] CPU.aluReg\[12\] _06906_ VGND VGND VPWR VPWR _06933_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14954__1032 clknet_1_0__leaf__02711_ VGND VGND VPWR VPWR net1064 sky130_fd_sc_hd__inv_2
X_11215_ _06316_ VGND VGND VPWR VPWR _01908_ sky130_fd_sc_hd__clkbuf_1
X_15176__1201 clknet_1_1__leaf__02748_ VGND VGND VPWR VPWR net1233 sky130_fd_sc_hd__inv_2
XFILLER_0_120_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12195_ CPU.aluReg\[30\] CPU.aluReg\[28\] _06871_ VGND VGND VPWR VPWR _06880_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11146_ CPU.registerFile\[8\]\[6\] _05723_ _06274_ VGND VGND VPWR VPWR _06280_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_50_Left_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15954_ CPU.registerFile\[9\]\[16\] _02802_ _03125_ VGND VGND VPWR VPWR _03437_ sky130_fd_sc_hd__o21a_1
X_11077_ net2508 _05723_ _06237_ VGND VGND VPWR VPWR _06243_ sky130_fd_sc_hd__mux2_1
X_14286__430 clknet_1_1__leaf__08462_ VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__inv_2
X_10028_ net1776 _05008_ _05607_ VGND VGND VPWR VPWR _05609_ sky130_fd_sc_hd__mux2_1
X_15885_ CPU.registerFile\[15\]\[14\] CPU.registerFile\[11\]\[14\] _02906_ VGND VGND
+ VPWR VPWR _03370_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17624_ net813 _01912_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[10\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_19_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17555_ net744 _01843_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_11979_ _06757_ VGND VGND VPWR VPWR _01582_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_868 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13718_ CPU.registerFile\[28\]\[24\] CPU.registerFile\[24\]\[24\] _07352_ VGND VGND
+ VPWR VPWR _08137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17486_ net675 _01774_ VGND VGND VPWR VPWR CPU.registerFile\[25\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16437_ CPU.registerFile\[1\]\[30\] _02867_ _03905_ _02895_ VGND VGND VPWR VPWR _03906_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13649_ _07519_ _08068_ _08069_ VGND VGND VPWR VPWR _08070_ sky130_fd_sc_hd__o21a_1
XFILLER_0_156_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14752__850 clknet_1_1__leaf__02691_ VGND VGND VPWR VPWR net882 sky130_fd_sc_hd__inv_2
X_16368_ CPU.registerFile\[30\]\[28\] CPU.registerFile\[26\]\[28\] _03247_ VGND VGND
+ VPWR VPWR _03839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18107_ net170 _02387_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15319_ _08403_ VGND VGND VPWR VPWR _02818_ sky130_fd_sc_hd__buf_4
XFILLER_0_30_908 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16512__180 clknet_1_0__leaf__03963_ VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__inv_2
X_16299_ CPU.registerFile\[5\]\[26\] CPU.registerFile\[4\]\[26\] _02806_ VGND VGND
+ VPWR VPWR _03772_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_113_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18038_ net1211 _02318_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_93_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09811_ net2112 _05230_ _05474_ VGND VGND VPWR VPWR _05477_ sky130_fd_sc_hd__mux2_1
X_09742_ _04478_ _04480_ VGND VGND VPWR VPWR _05431_ sky130_fd_sc_hd__nor2_1
X_09673_ _05361_ _05281_ _05364_ _05286_ VGND VGND VPWR VPWR _05365_ sky130_fd_sc_hd__o211a_1
X_08624_ _04248_ _04339_ _04340_ _04343_ VGND VGND VPWR VPWR _04344_ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ CPU.aluIn1\[6\] _04274_ VGND VGND VPWR VPWR _04275_ sky130_fd_sc_hd__and2_1
X_14835__925 clknet_1_1__leaf__02699_ VGND VGND VPWR VPWR net957 sky130_fd_sc_hd__inv_2
X_08486_ _04205_ VGND VGND VPWR VPWR _04206_ sky130_fd_sc_hd__buf_2
X_16576__49 clknet_1_0__leaf__03968_ VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__inv_2
XFILLER_0_147_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09107_ _04500_ _04292_ VGND VGND VPWR VPWR _04819_ sky130_fd_sc_hd__nand2_2
XFILLER_0_131_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09038_ _04357_ _04752_ _04671_ VGND VGND VPWR VPWR _04753_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_107_Left_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold360 CPU.registerFile\[28\]\[13\] VGND VGND VPWR VPWR net1601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 CPU.registerFile\[14\]\[18\] VGND VGND VPWR VPWR net1612 sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 CPU.PC\[12\] VGND VGND VPWR VPWR net1623 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold393 CPU.registerFile\[12\]\[12\] VGND VGND VPWR VPWR net1634 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ _06202_ VGND VGND VPWR VPWR _02009_ sky130_fd_sc_hd__clkbuf_1
X_14881__967 clknet_1_1__leaf__02703_ VGND VGND VPWR VPWR net999 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_144_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12951_ _04972_ VGND VGND VPWR VPWR _07392_ sky130_fd_sc_hd__buf_4
Xhold1060 CPU.registerFile\[31\]\[22\] VGND VGND VPWR VPWR net2301 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1071 CPU.registerFile\[21\]\[19\] VGND VGND VPWR VPWR net2312 sky130_fd_sc_hd__dlygate4sd3_1
X_11902_ net1657 _05681_ _06711_ VGND VGND VPWR VPWR _06717_ sky130_fd_sc_hd__mux2_1
X_15670_ CPU.registerFile\[8\]\[8\] _02763_ _03117_ _03160_ VGND VGND VPWR VPWR _03161_
+ sky130_fd_sc_hd__o211a_1
Xhold1082 CPU.registerFile\[21\]\[30\] VGND VGND VPWR VPWR net2323 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_200 _07841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_12882_ _07322_ _07323_ VGND VGND VPWR VPWR _07324_ sky130_fd_sc_hd__or2_1
Xhold1093 CPU.registerFile\[22\]\[30\] VGND VGND VPWR VPWR net2334 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_211 _07961_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_116_Left_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_222 clknet_1_0__leaf__02720_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_233 _02767_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11833_ _06680_ VGND VGND VPWR VPWR _01651_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_64_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_244 _03072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_255 _05045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_266 _05381_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17340_ net529 _01628_ VGND VGND VPWR VPWR CPU.registerFile\[10\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_277 _05551_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_288 _05727_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11764_ _04748_ net2520 _06639_ VGND VGND VPWR VPWR _06644_ sky130_fd_sc_hd__mux2_1
XANTENNA_299 _07320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13503_ CPU.registerFile\[21\]\[18\] _07502_ _07503_ CPU.registerFile\[17\]\[18\]
+ _07927_ VGND VGND VPWR VPWR _07928_ sky130_fd_sc_hd__o221a_1
X_10715_ _05522_ net1943 _06045_ VGND VGND VPWR VPWR _06051_ sky130_fd_sc_hd__mux2_1
X_17271_ clknet_leaf_13_clk _01559_ VGND VGND VPWR VPWR CPU.PC\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11695_ net2509 _06590_ _06600_ _06594_ VGND VGND VPWR VPWR _01708_ sky130_fd_sc_hd__o211a_1
XFILLER_0_138_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14474__600 clknet_1_1__leaf__02663_ VGND VGND VPWR VPWR net632 sky130_fd_sc_hd__inv_2
X_16222_ CPU.aluIn1\[23\] _02958_ _03680_ _03697_ _02995_ VGND VGND VPWR VPWR _02437_
+ sky130_fd_sc_hd__o221a_1
X_13434_ _07334_ _07851_ _07854_ _07861_ _07766_ VGND VGND VPWR VPWR _07862_ sky130_fd_sc_hd__o311a_1
XFILLER_0_82_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10646_ net1470 _05969_ VGND VGND VPWR VPWR _06008_ sky130_fd_sc_hd__or2_1
X_16153_ _08407_ _03607_ _03616_ _03630_ _07424_ VGND VGND VPWR VPWR _03631_ sky130_fd_sc_hd__a311o_2
Xrebuffer5 net1247 VGND VGND VPWR VPWR net1246 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13365_ CPU.registerFile\[31\]\[13\] _07276_ _07618_ CPU.registerFile\[27\]\[13\]
+ _07278_ VGND VGND VPWR VPWR _07795_ sky130_fd_sc_hd__o221a_1
XFILLER_0_106_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10577_ mapped_spi_flash.clk_div mapped_spi_flash.state\[3\] _05965_ VGND VGND VPWR
+ VPWR _05969_ sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_125_Left_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15104_ net1351 _07190_ VGND VGND VPWR VPWR _02739_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12316_ _06972_ VGND VGND VPWR VPWR _01425_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16084_ _08408_ _03554_ _03563_ _02993_ VGND VGND VPWR VPWR _03564_ sky130_fd_sc_hd__a31o_1
X_13296_ _07723_ _07724_ _07725_ _07727_ _07360_ VGND VGND VPWR VPWR _07728_ sky130_fd_sc_hd__a221o_1
XFILLER_0_139_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12247_ CPU.aluIn1\[17\] _06919_ _06894_ VGND VGND VPWR VPWR _06920_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12178_ net1291 _06865_ _06862_ _06867_ VGND VGND VPWR VPWR _01492_ sky130_fd_sc_hd__o211a_1
X_11129_ net2346 _05706_ _06263_ VGND VGND VPWR VPWR _06271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16986_ clknet_leaf_28_clk _01312_ VGND VGND VPWR VPWR CPU.rs2\[17\] sky130_fd_sc_hd__dfxtp_1
X_15158__1185 clknet_1_0__leaf__02746_ VGND VGND VPWR VPWR net1217 sky130_fd_sc_hd__inv_2
X_15937_ _02848_ _03416_ _03420_ _02843_ VGND VGND VPWR VPWR _03421_ sky130_fd_sc_hd__a211o_1
XFILLER_0_155_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_134_Left_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15868_ CPU.registerFile\[5\]\[13\] CPU.registerFile\[4\]\[13\] _03146_ VGND VGND
+ VPWR VPWR _03354_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_35_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17607_ net796 _01895_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[25\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_106_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15799_ CPU.registerFile\[5\]\[11\] CPU.registerFile\[4\]\[11\] _03146_ VGND VGND
+ VPWR VPWR _03287_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_106_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17538_ net727 _01826_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[20\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_156_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17469_ net658 _01757_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[24\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_921 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_126_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09725_ _04411_ _04300_ VGND VGND VPWR VPWR _05415_ sky130_fd_sc_hd__nand2_1
X_09656_ _04285_ _04211_ _04219_ CPU.aluReg\[4\] _05348_ VGND VGND VPWR VPWR _05349_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_2_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08607_ CPU.aluIn1\[13\] _04259_ VGND VGND VPWR VPWR _04327_ sky130_fd_sc_hd__and2_1
X_09587_ mapped_spi_ram.rcv_data\[14\] net18 _04618_ mapped_spi_flash.rcv_data\[14\]
+ VGND VGND VPWR VPWR _05282_ sky130_fd_sc_hd__a22o_2
X_14953__1031 clknet_1_1__leaf__02711_ VGND VGND VPWR VPWR net1063 sky130_fd_sc_hd__inv_2
X_14423__554 clknet_1_0__leaf__02658_ VGND VGND VPWR VPWR net586 sky130_fd_sc_hd__inv_2
X_08538_ CPU.aluIn1\[14\] _04257_ VGND VGND VPWR VPWR _04258_ sky130_fd_sc_hd__or2_1
X_15175__1200 clknet_1_1__leaf__02748_ VGND VGND VPWR VPWR net1232 sky130_fd_sc_hd__inv_2
XFILLER_0_64_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08469_ mapped_spi_ram.div_counter\[3\] mapped_spi_ram.div_counter\[2\] mapped_spi_ram.div_counter\[5\]
+ mapped_spi_ram.div_counter\[4\] VGND VGND VPWR VPWR _04191_ sky130_fd_sc_hd__nor4_1
XTAP_TAPCELL_ROW_42_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10500_ net1391 _05887_ _05856_ _05907_ VGND VGND VPWR VPWR _05908_ sky130_fd_sc_hd__a211o_1
XFILLER_0_18_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11480_ _06457_ VGND VGND VPWR VPWR _01784_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10431_ _05827_ VGND VGND VPWR VPWR _05851_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_21_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_154_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13150_ _07575_ _07585_ _07395_ VGND VGND VPWR VPWR _07586_ sky130_fd_sc_hd__o21a_1
X_10362_ _05539_ net2363 _05799_ VGND VGND VPWR VPWR _05803_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_749 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12101_ _06822_ VGND VGND VPWR VPWR _01524_ sky130_fd_sc_hd__clkbuf_1
X_10293_ _05539_ net2350 _05762_ VGND VGND VPWR VPWR _05766_ sky130_fd_sc_hd__mux2_1
X_13081_ _07272_ VGND VGND VPWR VPWR _07519_ sky130_fd_sc_hd__buf_4
XFILLER_0_103_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12032_ _04714_ net2211 _06783_ VGND VGND VPWR VPWR _06786_ sky130_fd_sc_hd__mux2_1
Xhold190 per_uart.uart0.enable16_counter\[14\] VGND VGND VPWR VPWR net1431 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16840_ _07195_ _03974_ VGND VGND VPWR VPWR _04137_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_70_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16771_ _04081_ _04085_ _04015_ VGND VGND VPWR VPWR _02598_ sky130_fd_sc_hd__a21oi_1
X_15722_ CPU.registerFile\[25\]\[9\] CPU.registerFile\[29\]\[9\] _02851_ VGND VGND
+ VPWR VPWR _03212_ sky130_fd_sc_hd__mux2_1
X_12934_ CPU.registerFile\[2\]\[2\] _07374_ VGND VGND VPWR VPWR _07375_ sky130_fd_sc_hd__or2_1
X_14506__629 clknet_1_1__leaf__02666_ VGND VGND VPWR VPWR net661 sky130_fd_sc_hd__inv_2
XFILLER_0_34_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15653_ CPU.registerFile\[2\]\[7\] _03143_ _02980_ CPU.registerFile\[3\]\[7\] _03144_
+ VGND VGND VPWR VPWR _03145_ sky130_fd_sc_hd__a221o_1
X_14244__417 clknet_1_1__leaf__08434_ VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__inv_2
X_12865_ _07126_ VGND VGND VPWR VPWR _07308_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_158_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_157_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11816_ _05402_ net1846 _06661_ VGND VGND VPWR VPWR _06671_ sky130_fd_sc_hd__mux2_1
X_18372_ net40 net31 VGND VGND VPWR VPWR mapped_spi_ram.div_counter\[4\] sky130_fd_sc_hd__dfxtp_1
X_15584_ _08410_ _03063_ _03077_ _02934_ VGND VGND VPWR VPWR _03078_ sky130_fd_sc_hd__o211a_1
X_12796_ _07238_ VGND VGND VPWR VPWR _07239_ sky130_fd_sc_hd__buf_4
XFILLER_0_56_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17323_ net512 _01611_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[19\] sky130_fd_sc_hd__dfxtp_1
X_14398__531 clknet_1_0__leaf__02656_ VGND VGND VPWR VPWR net563 sky130_fd_sc_hd__inv_2
XFILLER_0_141_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11747_ _06570_ _06633_ VGND VGND VPWR VPWR _06634_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17254_ net444 _01542_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_882 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11678_ net1478 _06590_ _06591_ _06581_ VGND VGND VPWR VPWR _01716_ sky130_fd_sc_hd__o211a_1
X_16205_ CPU.registerFile\[14\]\[23\] CPU.registerFile\[10\]\[23\] _02881_ VGND VGND
+ VPWR VPWR _03681_ sky130_fd_sc_hd__mux2_1
X_15074__1139 clknet_1_1__leaf__02723_ VGND VGND VPWR VPWR net1171 sky130_fd_sc_hd__inv_2
X_13417_ CPU.registerFile\[5\]\[15\] CPU.registerFile\[4\]\[15\] net14 VGND VGND VPWR
+ VPWR _07845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17185_ clknet_leaf_26_clk _01473_ VGND VGND VPWR VPWR CPU.Jimm\[15\] sky130_fd_sc_hd__dfxtp_1
X_10629_ mapped_spi_flash.rcv_data\[9\] _05994_ VGND VGND VPWR VPWR _05999_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16136_ CPU.registerFile\[25\]\[21\] _03280_ _02940_ VGND VGND VPWR VPWR _03614_
+ sky130_fd_sc_hd__o21a_1
X_13348_ CPU.registerFile\[6\]\[13\] CPU.registerFile\[7\]\[13\] _07263_ VGND VGND
+ VPWR VPWR _07778_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16067_ CPU.registerFile\[14\]\[19\] _02889_ VGND VGND VPWR VPWR _03547_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13279_ CPU.registerFile\[3\]\[11\] _07373_ _07710_ _07376_ VGND VGND VPWR VPWR _07711_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_90_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14864__951 clknet_1_0__leaf__02702_ VGND VGND VPWR VPWR net983 sky130_fd_sc_hd__inv_2
XFILLER_0_20_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_142_Left_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16969_ clknet_leaf_22_clk _01295_ VGND VGND VPWR VPWR CPU.mem_wdata\[0\] sky130_fd_sc_hd__dfxtp_2
X_09510_ _05208_ VGND VGND VPWR VPWR _05209_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_88_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09441_ _04435_ _04326_ VGND VGND VPWR VPWR _05143_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_88_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_121_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_121_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_760 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09372_ _04333_ _04256_ _05076_ VGND VGND VPWR VPWR _05077_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_821 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_151_Left_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_627 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_145_865 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_765 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_707 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16656__1 clknet_1_0__leaf__07220_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__inv_2
XFILLER_0_131_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09708_ _05393_ _05398_ _04708_ VGND VGND VPWR VPWR _05399_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_10980_ net1772 _05694_ _06190_ VGND VGND VPWR VPWR _06192_ sky130_fd_sc_hd__mux2_1
X_09639_ _05332_ VGND VGND VPWR VPWR _05333_ sky130_fd_sc_hd__buf_4
XFILLER_0_69_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12650_ _07150_ _07151_ VGND VGND VPWR VPWR _00018_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_26_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11601_ net1381 _06524_ _06538_ _06539_ VGND VGND VPWR VPWR _01741_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_139_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12581_ CPU.registerFile\[4\]\[5\] _05332_ _07107_ VGND VGND VPWR VPWR _07114_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_139_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11532_ _06482_ net1318 _06489_ _06492_ net1327 VGND VGND VPWR VPWR _01763_ sky130_fd_sc_hd__a32o_1
XFILLER_0_135_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15248__156 clknet_1_0__leaf__02755_ VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__inv_2
X_15157__1184 clknet_1_0__leaf__02746_ VGND VGND VPWR VPWR net1216 sky130_fd_sc_hd__inv_2
XFILLER_0_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11463_ _06448_ VGND VGND VPWR VPWR _01792_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_59_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13202_ net2384 _07358_ _07617_ _07636_ _05844_ VGND VGND VPWR VPWR _01303_ sky130_fd_sc_hd__o221a_1
XFILLER_0_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10414_ mapped_spi_flash.cmd_addr\[25\] _05825_ _05827_ mapped_spi_flash.cmd_addr\[26\]
+ VGND VGND VPWR VPWR _05839_ sky130_fd_sc_hd__a22o_1
X_11394_ _05518_ net2055 _06408_ VGND VGND VPWR VPWR _06412_ sky130_fd_sc_hd__mux2_1
X_13133_ CPU.registerFile\[21\]\[7\] _07362_ _07363_ CPU.registerFile\[17\]\[7\] _07568_
+ VGND VGND VPWR VPWR _07569_ sky130_fd_sc_hd__o221a_1
X_10345_ _05522_ net2396 _05788_ VGND VGND VPWR VPWR _05794_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14586__701 clknet_1_0__leaf__02674_ VGND VGND VPWR VPWR net733 sky130_fd_sc_hd__inv_2
XFILLER_0_103_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_72_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ _07235_ VGND VGND VPWR VPWR _07502_ sky130_fd_sc_hd__buf_4
X_17941_ net1130 _02225_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[21\] sky130_fd_sc_hd__dfxtp_1
X_10276_ _05522_ net1869 _05751_ VGND VGND VPWR VPWR _05757_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12015_ _06776_ VGND VGND VPWR VPWR _01565_ sky130_fd_sc_hd__clkbuf_1
X_17872_ net1061 _02156_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[30\] sky130_fd_sc_hd__dfxtp_1
X_16823_ _07195_ _07196_ _07197_ VGND VGND VPWR VPWR _04125_ sky130_fd_sc_hd__nor3_1
XFILLER_0_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16754_ _04032_ net1588 VGND VGND VPWR VPWR _04071_ sky130_fd_sc_hd__nand2_1
X_15705_ _02860_ VGND VGND VPWR VPWR _03195_ sky130_fd_sc_hd__buf_4
X_12917_ _07228_ VGND VGND VPWR VPWR _07358_ sky130_fd_sc_hd__buf_2
X_16685_ _04001_ _05319_ _03990_ VGND VGND VPWR VPWR _04013_ sky130_fd_sc_hd__a21o_1
X_13897_ CPU.registerFile\[14\]\[30\] CPU.registerFile\[10\]\[30\] _07480_ VGND VGND
+ VPWR VPWR _08310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_15636_ _03121_ _03127_ _02784_ VGND VGND VPWR VPWR _03128_ sky130_fd_sc_hd__a21o_1
X_12848_ _05337_ VGND VGND VPWR VPWR _07291_ sky130_fd_sc_hd__buf_4
XFILLER_0_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15567_ CPU.registerFile\[5\]\[5\] CPU.registerFile\[4\]\[5\] _02805_ VGND VGND VPWR
+ VPWR _03061_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_18355_ clknet_leaf_1_clk net1 VGND VGND VPWR VPWR per_uart.uart0.uart_rxd1 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17306_ net495 _01594_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_14518_ clknet_1_1__leaf__02664_ VGND VGND VPWR VPWR _02668_ sky130_fd_sc_hd__buf_1
XFILLER_0_124_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15498_ _02935_ _02985_ _02992_ _02993_ VGND VGND VPWR VPWR _02994_ sky130_fd_sc_hd__a31o_1
X_18286_ net119 _02566_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_154_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_17237_ net427 _01525_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_835 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_671 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold904 CPU.registerFile\[27\]\[23\] VGND VGND VPWR VPWR net2145 sky130_fd_sc_hd__dlygate4sd3_1
X_17168_ clknet_leaf_25_clk _01456_ VGND VGND VPWR VPWR CPU.mem_wmask\[0\] sky130_fd_sc_hd__dfxtp_1
Xhold915 CPU.registerFile\[8\]\[18\] VGND VGND VPWR VPWR net2156 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold926 CPU.registerFile\[10\]\[18\] VGND VGND VPWR VPWR net2167 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__08433_ _08433_ VGND VGND VPWR VPWR clknet_0__08433_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_51_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16119_ _08408_ _03588_ _03597_ _02993_ VGND VGND VPWR VPWR _03598_ sky130_fd_sc_hd__a31o_1
Xhold937 CPU.registerFile\[22\]\[23\] VGND VGND VPWR VPWR net2178 sky130_fd_sc_hd__dlygate4sd3_1
Xhold948 CPU.registerFile\[1\]\[19\] VGND VGND VPWR VPWR net2189 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09990_ _05545_ net2487 _05581_ VGND VGND VPWR VPWR _05588_ sky130_fd_sc_hd__mux2_1
X_17099_ net357 _01421_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[29\] sky130_fd_sc_hd__dfxtp_1
Xhold959 CPU.registerFile\[28\]\[6\] VGND VGND VPWR VPWR net2200 sky130_fd_sc_hd__dlygate4sd3_1
X_14452__580 clknet_1_0__leaf__02661_ VGND VGND VPWR VPWR net612 sky130_fd_sc_hd__inv_2
X_14952__1030 clknet_1_0__leaf__02711_ VGND VGND VPWR VPWR net1062 sky130_fd_sc_hd__inv_2
Xclkbuf_0__08364_ _08364_ VGND VGND VPWR VPWR clknet_0__08364_ sky130_fd_sc_hd__clkbuf_16
X_08941_ CPU.Bimm\[11\] VGND VGND VPWR VPWR _04661_ sky130_fd_sc_hd__buf_4
Xclkbuf_1_1__f__02688_ clknet_0__02688_ VGND VGND VPWR VPWR clknet_1_1__leaf__02688_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_4_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08872_ _04575_ _04590_ _04591_ _04586_ CPU.PC\[20\] VGND VGND VPWR VPWR _04592_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_126_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09424_ _04924_ _05126_ VGND VGND VPWR VPWR _05127_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09355_ _05057_ _05058_ _05060_ _04773_ VGND VGND VPWR VPWR _05061_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_23_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09286_ _04344_ _04994_ VGND VGND VPWR VPWR _04995_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14535__655 clknet_1_0__leaf__02669_ VGND VGND VPWR VPWR net687 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_134_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_10130_ net1556 _05359_ _05655_ VGND VGND VPWR VPWR _05663_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10061_ net2019 _05359_ _05618_ VGND VGND VPWR VPWR _05626_ sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f__03964_ clknet_0__03964_ VGND VGND VPWR VPWR clknet_1_0__leaf__03964_
+ sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_50_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13820_ CPU.registerFile\[8\]\[28\] CPU.registerFile\[12\]\[28\] _07233_ VGND VGND
+ VPWR VPWR _08235_ sky130_fd_sc_hd__mux2_1
X_15073__1138 clknet_1_1__leaf__02723_ VGND VGND VPWR VPWR net1170 sky130_fd_sc_hd__inv_2
XFILLER_0_98_844 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13751_ _07258_ _08166_ _08168_ _04987_ VGND VGND VPWR VPWR _08169_ sky130_fd_sc_hd__o211a_1
X_14581__697 clknet_1_1__leaf__02673_ VGND VGND VPWR VPWR net729 sky130_fd_sc_hd__inv_2
X_10963_ net1594 _05677_ _06179_ VGND VGND VPWR VPWR _06183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12702_ net1464 _07183_ VGND VGND VPWR VPWR _07184_ sky130_fd_sc_hd__or2_1
X_16470_ CPU.registerFile\[16\]\[31\] CPU.registerFile\[18\]\[31\] _05441_ VGND VGND
+ VPWR VPWR _03938_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13682_ CPU.registerFile\[1\]\[23\] _07387_ _08101_ _07379_ VGND VGND VPWR VPWR _08102_
+ sky130_fd_sc_hd__a211o_1
X_10894_ _06146_ VGND VGND VPWR VPWR _02059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_15421_ _02760_ VGND VGND VPWR VPWR _02918_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_155_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12633_ _07140_ net1356 VGND VGND VPWR VPWR _00042_ sky130_fd_sc_hd__nor2_1
XFILLER_0_155_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18140_ clknet_leaf_19_clk _02420_ VGND VGND VPWR VPWR CPU.aluIn1\[6\] sky130_fd_sc_hd__dfxtp_2
X_15352_ CPU.registerFile\[15\]\[1\] CPU.registerFile\[11\]\[1\] _02849_ VGND VGND
+ VPWR VPWR _02850_ sky130_fd_sc_hd__mux2_1
X_12564_ CPU.registerFile\[4\]\[13\] _05149_ _07096_ VGND VGND VPWR VPWR _07105_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11515_ _06478_ _06479_ _05855_ VGND VGND VPWR VPWR _01771_ sky130_fd_sc_hd__o21ai_1
X_18071_ net134 _02351_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_15283_ _05093_ VGND VGND VPWR VPWR _02782_ sky130_fd_sc_hd__clkbuf_4
X_12495_ _07068_ VGND VGND VPWR VPWR _01342_ sky130_fd_sc_hd__clkbuf_1
X_17022_ net280 _01344_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11446_ _06439_ VGND VGND VPWR VPWR _01800_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0__02711_ _02711_ VGND VGND VPWR VPWR clknet_0__02711_ sky130_fd_sc_hd__clkbuf_16
X_14165_ _08419_ VGND VGND VPWR VPWR _01483_ sky130_fd_sc_hd__clkbuf_1
X_11377_ _05501_ net1889 _06397_ VGND VGND VPWR VPWR _06403_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_150_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13116_ _07519_ _07551_ _07552_ VGND VGND VPWR VPWR _07553_ sky130_fd_sc_hd__o21a_1
X_10328_ _05505_ net2215 _05777_ VGND VGND VPWR VPWR _05785_ sky130_fd_sc_hd__mux2_1
X_14096_ _07128_ _08375_ VGND VGND VPWR VPWR _01458_ sky130_fd_sc_hd__nor2_1
XFILLER_0_147_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13047_ _07474_ _07479_ _07485_ VGND VGND VPWR VPWR _07486_ sky130_fd_sc_hd__or3_1
X_17924_ net1113 _02208_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[4\] sky130_fd_sc_hd__dfxtp_1
X_10259_ _05505_ net2121 _05740_ VGND VGND VPWR VPWR _05748_ sky130_fd_sc_hd__mux2_1
X_17855_ net1044 _02139_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[13\] sky130_fd_sc_hd__dfxtp_1
X_16806_ _04112_ _07200_ _07202_ _04113_ _06482_ VGND VGND VPWR VPWR _02605_ sky130_fd_sc_hd__o221ai_1
X_17786_ net975 _02070_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_844 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16737_ _04027_ _04039_ _05136_ VGND VGND VPWR VPWR _04057_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_85_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16668_ _03991_ net1562 VGND VGND VPWR VPWR _03998_ sky130_fd_sc_hd__nand2_1
XFILLER_0_158_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_146_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15619_ _02827_ _03110_ _03111_ VGND VGND VPWR VPWR _03112_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_45_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_16599_ clknet_1_0__leaf__07219_ VGND VGND VPWR VPWR _03971_ sky130_fd_sc_hd__buf_1
X_09140_ CPU.PC\[12\] _04851_ VGND VGND VPWR VPWR _04852_ sky130_fd_sc_hd__and2_1
X_18338_ clknet_leaf_2_clk _02618_ VGND VGND VPWR VPWR per_uart.rx_data\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09071_ _04709_ VGND VGND VPWR VPWR _04784_ sky130_fd_sc_hd__buf_4
X_18269_ clknet_leaf_1_clk _02549_ VGND VGND VPWR VPWR per_uart.uart0.rxd_reg\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold701 CPU.registerFile\[3\]\[13\] VGND VGND VPWR VPWR net1942 sky130_fd_sc_hd__dlygate4sd3_1
Xhold712 CPU.registerFile\[15\]\[23\] VGND VGND VPWR VPWR net1953 sky130_fd_sc_hd__dlygate4sd3_1
Xhold723 CPU.registerFile\[21\]\[4\] VGND VGND VPWR VPWR net1964 sky130_fd_sc_hd__dlygate4sd3_1
Xhold734 CPU.registerFile\[3\]\[19\] VGND VGND VPWR VPWR net1975 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold745 CPU.registerFile\[13\]\[12\] VGND VGND VPWR VPWR net1986 sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 CPU.registerFile\[27\]\[22\] VGND VGND VPWR VPWR net1997 sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 CPU.registerFile\[26\]\[2\] VGND VGND VPWR VPWR net2008 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold778 CPU.registerFile\[17\]\[4\] VGND VGND VPWR VPWR net2019 sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ _05528_ net1864 _05570_ VGND VGND VPWR VPWR _05579_ sky130_fd_sc_hd__mux2_1
Xhold789 CPU.registerFile\[29\]\[19\] VGND VGND VPWR VPWR net2030 sky130_fd_sc_hd__dlygate4sd3_1
X_08924_ _04635_ _04631_ _04641_ VGND VGND VPWR VPWR _04644_ sky130_fd_sc_hd__and3b_2
X_08855_ _04574_ _04571_ VGND VGND VPWR VPWR _04575_ sky130_fd_sc_hd__or2_4
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15156__1183 clknet_1_1__leaf__02746_ VGND VGND VPWR VPWR net1215 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f__02700_ clknet_0__02700_ VGND VGND VPWR VPWR clknet_1_0__leaf__02700_
+ sky130_fd_sc_hd__clkbuf_16
X_08786_ _04505_ CPU.state\[2\] CPU.state\[3\] VGND VGND VPWR VPWR _04506_ sky130_fd_sc_hd__or3_4
XFILLER_0_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09407_ _05110_ VGND VGND VPWR VPWR _02565_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09338_ _05040_ _05030_ _05031_ _05044_ VGND VGND VPWR VPWR _05045_ sky130_fd_sc_hd__or4b_4
XFILLER_0_35_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_893 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09269_ CPU.Iimm\[1\] _04812_ VGND VGND VPWR VPWR _04979_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11300_ _05493_ net2122 _06360_ VGND VGND VPWR VPWR _06362_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_12280_ _06945_ VGND VGND VPWR VPWR _01434_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_11231_ _06325_ VGND VGND VPWR VPWR _01901_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_11162_ _05487_ net1731 _06288_ VGND VGND VPWR VPWR _06289_ sky130_fd_sc_hd__mux2_1
X_10113_ CPU.registerFile\[18\]\[12\] _05170_ _05644_ VGND VGND VPWR VPWR _05654_
+ sky130_fd_sc_hd__mux2_1
X_11093_ _06251_ VGND VGND VPWR VPWR _06252_ sky130_fd_sc_hd__buf_4
X_15970_ CPU.registerFile\[1\]\[16\] _02939_ _03452_ _02894_ VGND VGND VPWR VPWR _03453_
+ sky130_fd_sc_hd__a22o_1
X_10044_ net2117 _05170_ _05607_ VGND VGND VPWR VPWR _05617_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold72 mapped_spi_ram.cmd_addr\[27\] VGND VGND VPWR VPWR net1313 sky130_fd_sc_hd__dlygate4sd3_1
X_17640_ net829 _01928_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[26\] sky130_fd_sc_hd__dfxtp_1
Xhold83 mapped_spi_flash.rcv_data\[20\] VGND VGND VPWR VPWR net1324 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 _06485_ VGND VGND VPWR VPWR net1335 sky130_fd_sc_hd__dlygate4sd3_1
X_14698__802 clknet_1_1__leaf__02685_ VGND VGND VPWR VPWR net834 sky130_fd_sc_hd__inv_2
X_13803_ _07646_ _08208_ _08211_ _08218_ VGND VGND VPWR VPWR _08219_ sky130_fd_sc_hd__a31o_1
X_17571_ net760 _01859_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_11995_ _05130_ net1689 _06758_ VGND VGND VPWR VPWR _06766_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_67_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13734_ CPU.registerFile\[1\]\[25\] _07619_ _08151_ _04939_ VGND VGND VPWR VPWR _08152_
+ sky130_fd_sc_hd__o22a_1
X_16522_ clknet_1_0__leaf__02749_ VGND VGND VPWR VPWR _03964_ sky130_fd_sc_hd__buf_1
X_10946_ _06173_ VGND VGND VPWR VPWR _02034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13665_ CPU.registerFile\[24\]\[23\] _07801_ _04987_ _08084_ VGND VGND VPWR VPWR
+ _08085_ sky130_fd_sc_hd__o211a_1
X_16453_ CPU.registerFile\[20\]\[30\] CPU.registerFile\[22\]\[30\] _05440_ VGND VGND
+ VPWR VPWR _03922_ sky130_fd_sc_hd__mux2_1
X_10877_ _06136_ VGND VGND VPWR VPWR _02066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_12616_ CPU.state\[1\] VGND VGND VPWR VPWR _07132_ sky130_fd_sc_hd__buf_2
X_15404_ _02895_ _02899_ _02900_ _02901_ VGND VGND VPWR VPWR _02902_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_80_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16384_ CPU.registerFile\[18\]\[28\] _02833_ _02836_ CPU.registerFile\[19\]\[28\]
+ _02910_ VGND VGND VPWR VPWR _03855_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_14_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13596_ _07228_ VGND VGND VPWR VPWR _08018_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_14_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15335_ _08394_ _05048_ VGND VGND VPWR VPWR _02834_ sky130_fd_sc_hd__nand2_2
X_18123_ net186 _02403_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[21\] sky130_fd_sc_hd__dfxtp_1
X_12547_ _07084_ VGND VGND VPWR VPWR _07096_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_81_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18054_ net1227 _02334_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[16\] sky130_fd_sc_hd__dfxtp_1
X_15266_ CPU.registerFile\[12\]\[0\] _05049_ VGND VGND VPWR VPWR _02765_ sky130_fd_sc_hd__or2_1
X_12478_ _07059_ VGND VGND VPWR VPWR _01350_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_3 CPU.mem_wdata\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_17005_ clknet_leaf_7_clk net1342 VGND VGND VPWR VPWR per_uart.uart0.enable16_counter\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_11429_ _05553_ net1654 _06396_ VGND VGND VPWR VPWR _06430_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15197_ clknet_1_1__leaf__02749_ VGND VGND VPWR VPWR _02751_ sky130_fd_sc_hd__buf_1
XFILLER_0_10_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14148_ _08409_ VGND VGND VPWR VPWR _01476_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_158_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17907_ net1096 _02191_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[25\] sky130_fd_sc_hd__dfxtp_1
X_08640_ _04357_ _04232_ _04359_ VGND VGND VPWR VPWR _04360_ sky130_fd_sc_hd__o21a_1
X_17838_ net1027 _02122_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[28\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer15 net1257 VGND VGND VPWR VPWR net1256 sky130_fd_sc_hd__dlygate4sd1_1
X_14564__681 clknet_1_1__leaf__02672_ VGND VGND VPWR VPWR net713 sky130_fd_sc_hd__inv_2
Xrebuffer26 net1268 VGND VGND VPWR VPWR net1267 sky130_fd_sc_hd__clkbuf_2
X_08571_ CPU.instr\[6\] VGND VGND VPWR VPWR _04291_ sky130_fd_sc_hd__buf_2
Xrebuffer37 _04538_ VGND VGND VPWR VPWR net1278 sky130_fd_sc_hd__dlygate4sd1_1
X_17769_ net958 _02053_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[23\] sky130_fd_sc_hd__dfxtp_1
Xrebuffer48 _04203_ VGND VGND VPWR VPWR net1295 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_09123_ _04833_ _04834_ VGND VGND VPWR VPWR _04835_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09054_ _04677_ VGND VGND VPWR VPWR _04768_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15072__1137 clknet_1_1__leaf__02723_ VGND VGND VPWR VPWR net1169 sky130_fd_sc_hd__inv_2
Xhold520 CPU.registerFile\[28\]\[26\] VGND VGND VPWR VPWR net1761 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold531 CPU.registerFile\[6\]\[20\] VGND VGND VPWR VPWR net1772 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold542 CPU.registerFile\[3\]\[3\] VGND VGND VPWR VPWR net1783 sky130_fd_sc_hd__dlygate4sd3_1
Xhold553 CPU.registerFile\[26\]\[6\] VGND VGND VPWR VPWR net1794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 CPU.registerFile\[20\]\[30\] VGND VGND VPWR VPWR net1805 sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 CPU.registerFile\[5\]\[2\] VGND VGND VPWR VPWR net1816 sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 CPU.registerFile\[3\]\[12\] VGND VGND VPWR VPWR net1827 sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 CPU.registerFile\[14\]\[19\] VGND VGND VPWR VPWR net1838 sky130_fd_sc_hd__dlygate4sd3_1
X_09956_ _05558_ VGND VGND VPWR VPWR _05570_ sky130_fd_sc_hd__buf_4
X_14647__756 clknet_1_1__leaf__02680_ VGND VGND VPWR VPWR net788 sky130_fd_sc_hd__inv_2
X_08907_ _04530_ _04626_ VGND VGND VPWR VPWR _04627_ sky130_fd_sc_hd__nand2_1
X_09887_ _05129_ VGND VGND VPWR VPWR _05526_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_129_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1220 CPU.registerFile\[19\]\[13\] VGND VGND VPWR VPWR net2461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1231 CPU.registerFile\[25\]\[2\] VGND VGND VPWR VPWR net2472 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1242 CPU.registerFile\[4\]\[26\] VGND VGND VPWR VPWR net2483 sky130_fd_sc_hd__dlygate4sd3_1
X_08838_ _04555_ _04554_ _04553_ _04556_ _04557_ VGND VGND VPWR VPWR _04558_ sky130_fd_sc_hd__o311ai_4
Xhold1253 CPU.registerFile\[21\]\[1\] VGND VGND VPWR VPWR net2494 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_142_Right_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1264 mapped_spi_flash.rcv_data\[8\] VGND VGND VPWR VPWR net2505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1275 CPU.registerFile\[20\]\[9\] VGND VGND VPWR VPWR net2516 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1286 CPU.aluReg\[27\] VGND VGND VPWR VPWR net2527 sky130_fd_sc_hd__dlygate4sd3_1
X_08769_ _04488_ VGND VGND VPWR VPWR _04489_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_404 _03138_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1297 mapped_spi_flash.cmd_addr\[25\] VGND VGND VPWR VPWR net2538 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_415 _05333_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_142_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ _05539_ net1773 _06092_ VGND VGND VPWR VPWR _06096_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_49_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _06652_ VGND VGND VPWR VPWR _01676_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10731_ _06059_ VGND VGND VPWR VPWR _02135_ sky130_fd_sc_hd__clkbuf_1
X_13450_ _07380_ _07872_ _07876_ _07584_ VGND VGND VPWR VPWR _07877_ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10662_ mapped_spi_flash.rcv_bitcount\[4\] _05964_ mapped_spi_flash.state\[3\] VGND
+ VGND VPWR VPWR _06020_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_62_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12401_ _04762_ net2161 _07013_ VGND VGND VPWR VPWR _07019_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14693__798 clknet_1_1__leaf__02684_ VGND VGND VPWR VPWR net830 sky130_fd_sc_hd__inv_2
XFILLER_0_24_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_14021__300 clknet_1_1__leaf__08362_ VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__inv_2
X_13381_ CPU.registerFile\[18\]\[14\] CPU.registerFile\[22\]\[14\] _07457_ VGND VGND
+ VPWR VPWR _07810_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_790 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_872 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_10593_ net1475 _05970_ VGND VGND VPWR VPWR _05978_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14392__526 clknet_1_0__leaf__02655_ VGND VGND VPWR VPWR net558 sky130_fd_sc_hd__inv_2
XFILLER_0_51_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12332_ _06982_ VGND VGND VPWR VPWR _01419_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12263_ _06932_ VGND VGND VPWR VPWR _01438_ sky130_fd_sc_hd__clkbuf_1
Xoutput5 net5 VGND VGND VPWR VPWR LEDS sky130_fd_sc_hd__clkbuf_4
X_11214_ _05543_ net2274 _06310_ VGND VGND VPWR VPWR _06316_ sky130_fd_sc_hd__mux2_1
X_12194_ _06879_ VGND VGND VPWR VPWR _01454_ sky130_fd_sc_hd__clkbuf_1
X_11145_ _06279_ VGND VGND VPWR VPWR _01941_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15953_ CPU.registerFile\[13\]\[16\] _03123_ VGND VGND VPWR VPWR _03436_ sky130_fd_sc_hd__or2_1
X_11076_ _06242_ VGND VGND VPWR VPWR _01973_ sky130_fd_sc_hd__clkbuf_1
X_10027_ _05608_ VGND VGND VPWR VPWR _02403_ sky130_fd_sc_hd__clkbuf_1
X_15884_ _02759_ _03366_ _03368_ _03019_ VGND VGND VPWR VPWR _03369_ sky130_fd_sc_hd__a211o_1
X_17623_ net812 _01911_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_28_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_19_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17554_ net743 _01842_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_11978_ _04958_ net2066 _06747_ VGND VGND VPWR VPWR _06757_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10929_ _06164_ VGND VGND VPWR VPWR _02042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_817 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13717_ CPU.registerFile\[29\]\[24\] _07347_ _07348_ CPU.registerFile\[25\]\[24\]
+ _07300_ VGND VGND VPWR VPWR _08136_ sky130_fd_sc_hd__o221a_1
X_17485_ net674 _01773_ VGND VGND VPWR VPWR mapped_spi_ram.rbusy sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16436_ CPU.registerFile\[5\]\[30\] CPU.registerFile\[4\]\[30\] _02806_ VGND VGND
+ VPWR VPWR _03905_ sky130_fd_sc_hd__mux2_1
X_13648_ CPU.registerFile\[13\]\[22\] _07361_ _07521_ CPU.registerFile\[9\]\[22\]
+ _07554_ VGND VGND VPWR VPWR _08069_ sky130_fd_sc_hd__o221a_1
XFILLER_0_27_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_13579_ CPU.registerFile\[15\]\[20\] _07236_ _07277_ CPU.registerFile\[11\]\[20\]
+ _07820_ VGND VGND VPWR VPWR _08002_ sky130_fd_sc_hd__o221a_1
X_16367_ _03833_ _03837_ _08410_ VGND VGND VPWR VPWR _03838_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_883 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_143_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18106_ net169 _02386_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15318_ CPU.registerFile\[1\]\[0\] _02814_ _02815_ _02816_ VGND VGND VPWR VPWR _02817_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16298_ _08397_ _03766_ _03770_ _02903_ VGND VGND VPWR VPWR _03771_ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15155__1182 clknet_1_0__leaf__02746_ VGND VGND VPWR VPWR net1214 sky130_fd_sc_hd__inv_2
XFILLER_0_78_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18037_ net1210 _02317_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_55 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_93_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09810_ _05476_ VGND VGND VPWR VPWR _02520_ sky130_fd_sc_hd__clkbuf_1
X_14369__506 clknet_1_1__leaf__02652_ VGND VGND VPWR VPWR net538 sky130_fd_sc_hd__inv_2
X_09741_ _05417_ _04716_ _05428_ _05429_ VGND VGND VPWR VPWR _05430_ sky130_fd_sc_hd__a31o_1
X_09672_ _04625_ _05173_ _05277_ _05363_ VGND VGND VPWR VPWR _05364_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_97_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08623_ _04341_ _04342_ VGND VGND VPWR VPWR _04343_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_19_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_38_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_08554_ CPU.mem_wdata\[6\] CPU.Bimm\[6\] _04203_ VGND VGND VPWR VPWR _04274_ sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_124_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08485_ _04204_ VGND VGND VPWR VPWR _04205_ sky130_fd_sc_hd__buf_2
XFILLER_0_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09106_ _04817_ VGND VGND VPWR VPWR _04818_ sky130_fd_sc_hd__buf_2
XFILLER_0_134_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_131_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_09037_ _04356_ _04234_ _04354_ VGND VGND VPWR VPWR _04752_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold350 per_uart.uart0.rxd_reg\[5\] VGND VGND VPWR VPWR net1591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 CPU.registerFile\[4\]\[2\] VGND VGND VPWR VPWR net1602 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold372 CPU.registerFile\[16\]\[27\] VGND VGND VPWR VPWR net1613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 CPU.registerFile\[14\]\[20\] VGND VGND VPWR VPWR net1624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 mapped_spi_ram.rcv_data\[3\] VGND VGND VPWR VPWR net1635 sky130_fd_sc_hd__dlygate4sd3_1
X_09939_ _05561_ VGND VGND VPWR VPWR _02476_ sky130_fd_sc_hd__clkbuf_1
X_16639__84 clknet_1_0__leaf__03988_ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_144_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12950_ CPU.registerFile\[1\]\[2\] _07387_ _07390_ _07231_ VGND VGND VPWR VPWR _07391_
+ sky130_fd_sc_hd__a211o_1
Xhold1050 CPU.registerFile\[3\]\[24\] VGND VGND VPWR VPWR net2291 sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ _06716_ VGND VGND VPWR VPWR _01619_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1061 CPU.registerFile\[21\]\[20\] VGND VGND VPWR VPWR net2302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1072 CPU.cycles\[10\] VGND VGND VPWR VPWR net2313 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1083 CPU.registerFile\[15\]\[13\] VGND VGND VPWR VPWR net2324 sky130_fd_sc_hd__dlygate4sd3_1
X_16654__98 clknet_1_1__leaf__03989_ VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__inv_2
X_12881_ CPU.registerFile\[18\]\[1\] CPU.registerFile\[22\]\[1\] _05283_ VGND VGND
+ VPWR VPWR _07323_ sky130_fd_sc_hd__mux2_1
Xhold1094 CPU.registerFile\[22\]\[29\] VGND VGND VPWR VPWR net2335 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_201 _07841_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_212 _07984_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_223 clknet_1_0__leaf__02720_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_11832_ net1862 _05679_ _06675_ VGND VGND VPWR VPWR _06680_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_16_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_234 _02775_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_245 _03091_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_256 _05045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_267 _05381_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_14551_ clknet_1_0__leaf__02664_ VGND VGND VPWR VPWR _02671_ sky130_fd_sc_hd__buf_1
X_11763_ _06643_ VGND VGND VPWR VPWR _01684_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_278 _05551_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_289 _05727_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10714_ _06050_ VGND VGND VPWR VPWR _02143_ sky130_fd_sc_hd__clkbuf_1
X_13502_ _07245_ _07926_ VGND VGND VPWR VPWR _07927_ sky130_fd_sc_hd__or2_1
X_17270_ net460 _01558_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11694_ mapped_spi_ram.rcv_data\[13\] _06588_ VGND VGND VPWR VPWR _06600_ sky130_fd_sc_hd__or2_1
X_14400__533 clknet_1_0__leaf__02656_ VGND VGND VPWR VPWR net565 sky130_fd_sc_hd__inv_2
XFILLER_0_36_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_16221_ _08408_ _03688_ _03696_ _02993_ VGND VGND VPWR VPWR _03697_ sky130_fd_sc_hd__a31o_1
X_13433_ _07555_ _07857_ _07858_ _07860_ _07302_ VGND VGND VPWR VPWR _07861_ sky130_fd_sc_hd__a221o_2
X_10645_ net1470 _05996_ _06007_ _06006_ VGND VGND VPWR VPWR _02168_ sky130_fd_sc_hd__o211a_1
XFILLER_0_24_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16152_ _02936_ _03622_ _03629_ _02843_ VGND VGND VPWR VPWR _03630_ sky130_fd_sc_hd__o211a_1
X_13364_ CPU.registerFile\[29\]\[13\] _07289_ _07290_ CPU.registerFile\[25\]\[13\]
+ _07793_ VGND VGND VPWR VPWR _07794_ sky130_fd_sc_hd__o221a_1
XFILLER_0_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer6 net1248 VGND VGND VPWR VPWR net1247 sky130_fd_sc_hd__clkbuf_2
X_10576_ _05967_ VGND VGND VPWR VPWR _05968_ sky130_fd_sc_hd__buf_2
XFILLER_0_24_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15103_ _07190_ net1446 _02727_ VGND VGND VPWR VPWR _02281_ sky130_fd_sc_hd__a21oi_1
X_12315_ CPU.aluReg\[1\] _06971_ _06861_ VGND VGND VPWR VPWR _06972_ sky130_fd_sc_hd__mux2_1
X_16083_ _03558_ _03562_ _02810_ VGND VGND VPWR VPWR _03563_ sky130_fd_sc_hd__a21o_1
X_13295_ _07398_ _07726_ VGND VGND VPWR VPWR _07727_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12246_ CPU.aluReg\[18\] CPU.aluReg\[16\] _06906_ VGND VGND VPWR VPWR _06919_ sky130_fd_sc_hd__mux2_1
XFILLER_0_139_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12177_ net2374 _06866_ VGND VGND VPWR VPWR _06867_ sky130_fd_sc_hd__xor2_1
X_11128_ _06270_ VGND VGND VPWR VPWR _01949_ sky130_fd_sc_hd__clkbuf_1
X_16985_ clknet_leaf_29_clk _01311_ VGND VGND VPWR VPWR CPU.rs2\[16\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11059_ _06233_ VGND VGND VPWR VPWR _01981_ sky130_fd_sc_hd__clkbuf_1
X_15936_ _03015_ _03417_ _03419_ _03019_ VGND VGND VPWR VPWR _03420_ sky130_fd_sc_hd__o211a_1
X_15867_ CPU.registerFile\[2\]\[13\] _03143_ _02980_ CPU.registerFile\[3\]\[13\] _03144_
+ VGND VGND VPWR VPWR _03353_ sky130_fd_sc_hd__a221o_1
X_15071__1136 clknet_1_1__leaf__02723_ VGND VGND VPWR VPWR net1168 sky130_fd_sc_hd__inv_2
XFILLER_0_154_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17606_ net795 _01894_ VGND VGND VPWR VPWR CPU.registerFile\[9\]\[24\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_35_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14818_ clknet_1_0__leaf__02697_ VGND VGND VPWR VPWR _02698_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_106_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15798_ CPU.registerFile\[2\]\[11\] _03143_ _02980_ CPU.registerFile\[3\]\[11\] _03144_
+ VGND VGND VPWR VPWR _03286_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_106_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17537_ net726 _01825_ VGND VGND VPWR VPWR CPU.registerFile\[24\]\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_17468_ net657 _01756_ VGND VGND VPWR VPWR mapped_spi_ram.cmd_addr\[23\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_14676__782 clknet_1_1__leaf__02683_ VGND VGND VPWR VPWR net814 sky130_fd_sc_hd__inv_2
X_16419_ CPU.registerFile\[27\]\[29\] _02928_ _02923_ VGND VGND VPWR VPWR _03889_
+ sky130_fd_sc_hd__o21a_1
X_14375__510 clknet_1_0__leaf__02654_ VGND VGND VPWR VPWR net542 sky130_fd_sc_hd__inv_2
X_17399_ net588 _01687_ VGND VGND VPWR VPWR CPU.registerFile\[13\]\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16581__53 clknet_1_0__leaf__03969_ VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__inv_2
XFILLER_0_15_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_113_933 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_8_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_8
X_14074__348 clknet_1_0__leaf__08367_ VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__inv_2
XFILLER_0_59_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14841__930 clknet_1_1__leaf__02700_ VGND VGND VPWR VPWR net962 sky130_fd_sc_hd__inv_2
X_09724_ CPU.cycles\[1\] _04989_ _05290_ CPU.PC\[1\] _05413_ VGND VGND VPWR VPWR _05414_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_126_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09655_ _04308_ _04683_ VGND VGND VPWR VPWR _05348_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_2_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_08606_ _04324_ _04262_ _04325_ VGND VGND VPWR VPWR _04326_ sky130_fd_sc_hd__a21o_1
XFILLER_0_145_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09586_ _04208_ _04624_ _05280_ VGND VGND VPWR VPWR _05281_ sky130_fd_sc_hd__o21ai_2
X_14759__857 clknet_1_1__leaf__02691_ VGND VGND VPWR VPWR net889 sky130_fd_sc_hd__inv_2
X_08537_ CPU.rs2\[14\] _04200_ _04205_ VGND VGND VPWR VPWR _04257_ sky130_fd_sc_hd__a21o_1
XFILLER_0_93_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16519__187 clknet_1_0__leaf__03963_ VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_42_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10430_ _05817_ VGND VGND VPWR VPWR _05850_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_154_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10361_ _05802_ VGND VGND VPWR VPWR _02248_ sky130_fd_sc_hd__clkbuf_1
X_12100_ _04714_ net2400 _06819_ VGND VGND VPWR VPWR _06822_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13080_ _07273_ _07516_ _07517_ VGND VGND VPWR VPWR _07518_ sky130_fd_sc_hd__o21a_1
X_10292_ _05765_ VGND VGND VPWR VPWR _02295_ sky130_fd_sc_hd__clkbuf_1
X_12031_ _06785_ VGND VGND VPWR VPWR _01557_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_57_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold180 CPU.cycles\[29\] VGND VGND VPWR VPWR net1421 sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 _02741_ VGND VGND VPWR VPWR net1432 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_16770_ _04050_ _04082_ _04083_ _04084_ VGND VGND VPWR VPWR _04085_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_70_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15721_ CPU.registerFile\[27\]\[9\] CPU.registerFile\[31\]\[9\] _02852_ VGND VGND
+ VPWR VPWR _03211_ sky130_fd_sc_hd__mux2_1
X_12933_ _05337_ VGND VGND VPWR VPWR _07374_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_15154__1181 clknet_1_1__leaf__02746_ VGND VGND VPWR VPWR net1213 sky130_fd_sc_hd__inv_2
X_15652_ _02779_ VGND VGND VPWR VPWR _03144_ sky130_fd_sc_hd__clkbuf_4
X_12864_ _07271_ _07280_ _07287_ _07303_ _07306_ VGND VGND VPWR VPWR _07307_ sky130_fd_sc_hd__o311a_1
X_11815_ _06670_ VGND VGND VPWR VPWR _01659_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18371_ net39 net30 VGND VGND VPWR VPWR mapped_spi_ram.div_counter\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_157_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_828 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12795_ _07237_ VGND VGND VPWR VPWR _07238_ sky130_fd_sc_hd__buf_2
XFILLER_0_139_841 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15583_ _02948_ _03071_ _03076_ VGND VGND VPWR VPWR _03077_ sky130_fd_sc_hd__or3_2
X_17322_ net511 _01610_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11746_ net2542 mapped_spi_ram.rcv_bitcount\[0\] net1349 VGND VGND VPWR VPWR _06633_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17253_ net443 _01541_ VGND VGND VPWR VPWR CPU.registerFile\[26\]\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_59 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11677_ net1448 _06588_ VGND VGND VPWR VPWR _06591_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_16204_ _02935_ _03679_ VGND VGND VPWR VPWR _03680_ sky130_fd_sc_hd__and2_1
X_13416_ _07842_ _07843_ _07476_ VGND VGND VPWR VPWR _07844_ sky130_fd_sc_hd__mux2_1
X_10628_ net2441 _05996_ _05998_ _05993_ VGND VGND VPWR VPWR _02176_ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_14396_ clknet_1_0__leaf__02653_ VGND VGND VPWR VPWR _02656_ sky130_fd_sc_hd__buf_1
X_17184_ clknet_leaf_14_clk _01472_ VGND VGND VPWR VPWR CPU.Jimm\[14\] sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_40_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_13347_ _07771_ _07776_ _07320_ VGND VGND VPWR VPWR _07777_ sky130_fd_sc_hd__mux2_1
X_16135_ CPU.registerFile\[29\]\[21\] _02918_ VGND VGND VPWR VPWR _03613_ sky130_fd_sc_hd__or2_1
X_10559_ net1452 _05943_ VGND VGND VPWR VPWR _05955_ sky130_fd_sc_hd__nand2_1
X_15225__135 clknet_1_1__leaf__02753_ VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__inv_2
XFILLER_0_121_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13278_ CPU.registerFile\[2\]\[11\] _07374_ VGND VGND VPWR VPWR _07710_ sky130_fd_sc_hd__or2_1
X_16066_ CPU.registerFile\[8\]\[19\] CPU.registerFile\[12\]\[19\] _03254_ VGND VGND
+ VPWR VPWR _03546_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_12229_ _06870_ VGND VGND VPWR VPWR _06906_ sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_90_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15017_ clknet_1_1__leaf__02708_ VGND VGND VPWR VPWR _02717_ sky130_fd_sc_hd__buf_1
X_16968_ net263 _01294_ VGND VGND VPWR VPWR CPU.registerFile\[4\]\[31\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_108_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15919_ CPU.registerFile\[11\]\[15\] _02861_ VGND VGND VPWR VPWR _03403_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16899_ CPU.mem_wdata\[0\] _04174_ _04175_ _04176_ VGND VGND VPWR VPWR _02635_ sky130_fd_sc_hd__o211a_1
X_09440_ _04260_ _04211_ _04681_ CPU.aluReg\[13\] _05141_ VGND VGND VPWR VPWR _05142_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_88_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16633__79 clknet_1_0__leaf__03971_ VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_121_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09371_ _04332_ _04330_ VGND VGND VPWR VPWR _05076_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_772 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_877 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_140_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09707_ net1294 _04489_ _05397_ _04679_ VGND VGND VPWR VPWR _05398_ sky130_fd_sc_hd__a22o_1
X_09638_ _05316_ _05325_ _05331_ VGND VGND VPWR VPWR _05332_ sky130_fd_sc_hd__or3b_4
X_14347__486 clknet_1_1__leaf__08467_ VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__inv_2
XFILLER_0_85_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09569_ _04800_ _05261_ _05264_ _04678_ VGND VGND VPWR VPWR _05265_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_26_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13985__268 clknet_1_0__leaf__08358_ VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__inv_2
X_11600_ _06515_ VGND VGND VPWR VPWR _06539_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_26_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12580_ _07113_ VGND VGND VPWR VPWR _01269_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_800 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_139_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_156_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_156_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_11531_ _06482_ net2541 _06489_ _06492_ net1318 VGND VGND VPWR VPWR _01764_ sky130_fd_sc_hd__a32o_1
XFILLER_0_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16545__20 clknet_1_0__leaf__03966_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__inv_2
X_11462_ _05518_ net2206 _06444_ VGND VGND VPWR VPWR _06448_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13201_ _07397_ _07627_ _07635_ _07424_ VGND VGND VPWR VPWR _07636_ sky130_fd_sc_hd__a31o_2
XTAP_TAPCELL_ROW_59_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10413_ _05838_ VGND VGND VPWR VPWR _02231_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_59_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_11393_ _06411_ VGND VGND VPWR VPWR _01825_ sky130_fd_sc_hd__clkbuf_1
X_16560__34 clknet_1_0__leaf__03967_ VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__inv_2
X_15070__1135 clknet_1_0__leaf__02723_ VGND VGND VPWR VPWR net1167 sky130_fd_sc_hd__inv_2
X_13132_ _07364_ _07567_ VGND VGND VPWR VPWR _07568_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_10344_ _05793_ VGND VGND VPWR VPWR _02256_ sky130_fd_sc_hd__clkbuf_1
X_14057__332 clknet_1_0__leaf__08366_ VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__inv_2
X_14512__634 clknet_1_0__leaf__02667_ VGND VGND VPWR VPWR net666 sky130_fd_sc_hd__inv_2
XFILLER_0_29_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17940_ net1129 _02224_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[20\] sky130_fd_sc_hd__dfxtp_1
X_13063_ CPU.registerFile\[23\]\[5\] _07325_ _07500_ CPU.registerFile\[19\]\[5\] _07327_
+ VGND VGND VPWR VPWR _07501_ sky130_fd_sc_hd__o221a_1
X_10275_ _05756_ VGND VGND VPWR VPWR _02303_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_72_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_14250__422 clknet_1_1__leaf__08435_ VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__inv_2
X_12014_ _05333_ net2173 _06769_ VGND VGND VPWR VPWR _06776_ sky130_fd_sc_hd__mux2_1
X_17871_ net1060 _02155_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[29\] sky130_fd_sc_hd__dfxtp_1
X_16822_ _04123_ _04122_ _04124_ _03632_ VGND VGND VPWR VPWR _02610_ sky130_fd_sc_hd__o211a_1
X_16753_ _04066_ _04070_ _05942_ VGND VGND VPWR VPWR _02595_ sky130_fd_sc_hd__o21a_1
X_13965_ clknet_1_1__leaf__07223_ VGND VGND VPWR VPWR _08357_ sky130_fd_sc_hd__buf_1
X_15704_ _03192_ _03193_ _02856_ VGND VGND VPWR VPWR _03194_ sky130_fd_sc_hd__mux2_1
X_12916_ CPU.mem_wdata\[1\] _07229_ _07357_ _07135_ VGND VGND VPWR VPWR _01296_ sky130_fd_sc_hd__o211a_1
X_16684_ _08379_ _05327_ _04006_ VGND VGND VPWR VPWR _04012_ sky130_fd_sc_hd__or3b_1
X_13896_ _08302_ _08308_ _07514_ VGND VGND VPWR VPWR _08309_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_103_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_15635_ _02771_ _03122_ _03124_ _03126_ _02782_ VGND VGND VPWR VPWR _03127_ sky130_fd_sc_hd__a221o_1
XFILLER_0_69_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_12847_ _07238_ VGND VGND VPWR VPWR _07290_ sky130_fd_sc_hd__buf_4
XFILLER_0_56_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_18354_ clknet_leaf_5_clk _02634_ VGND VGND VPWR VPWR per_uart.rx_avail sky130_fd_sc_hd__dfxtp_1
X_15566_ CPU.registerFile\[2\]\[5\] _02872_ _02980_ CPU.registerFile\[3\]\[5\] _02940_
+ VGND VGND VPWR VPWR _03060_ sky130_fd_sc_hd__a221o_1
XFILLER_0_127_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_139_682 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17305_ net494 _01593_ VGND VGND VPWR VPWR CPU.registerFile\[11\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18285_ net118 _02565_ VGND VGND VPWR VPWR CPU.registerFile\[16\]\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11729_ _06619_ net1310 VGND VGND VPWR VPWR _06621_ sky130_fd_sc_hd__and2b_1
XFILLER_0_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15497_ _07308_ VGND VGND VPWR VPWR _02993_ sky130_fd_sc_hd__buf_4
X_17236_ net426 _01524_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[29\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_142_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_141_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17167_ net391 _01455_ VGND VGND VPWR VPWR CPU.aluReg\[31\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_869 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold905 CPU.registerFile\[7\]\[7\] VGND VGND VPWR VPWR net2146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold916 CPU.registerFile\[17\]\[18\] VGND VGND VPWR VPWR net2157 sky130_fd_sc_hd__dlygate4sd3_1
Xhold927 CPU.registerFile\[15\]\[10\] VGND VGND VPWR VPWR net2168 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_0__08432_ _08432_ VGND VGND VPWR VPWR clknet_0__08432_ sky130_fd_sc_hd__clkbuf_16
X_16118_ _03592_ _03596_ _02810_ VGND VGND VPWR VPWR _03597_ sky130_fd_sc_hd__a21o_1
Xhold938 CPU.registerFile\[1\]\[1\] VGND VGND VPWR VPWR net2179 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17098_ net356 _01420_ VGND VGND VPWR VPWR CPU.registerFile\[29\]\[28\] sky130_fd_sc_hd__dfxtp_1
Xhold949 CPU.registerFile\[24\]\[15\] VGND VGND VPWR VPWR net2190 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f__02756_ clknet_0__02756_ VGND VGND VPWR VPWR clknet_1_1__leaf__02756_
+ sky130_fd_sc_hd__clkbuf_16
X_14788__883 clknet_1_1__leaf__02694_ VGND VGND VPWR VPWR net915 sky130_fd_sc_hd__inv_2
Xclkbuf_0__08363_ _08363_ VGND VGND VPWR VPWR clknet_0__08363_ sky130_fd_sc_hd__clkbuf_16
X_16049_ _08407_ _03506_ _03515_ _03529_ _07424_ VGND VGND VPWR VPWR _03530_ sky130_fd_sc_hd__a311o_2
X_08940_ CPU.Bimm\[1\] VGND VGND VPWR VPWR _04660_ sky130_fd_sc_hd__buf_4
XFILLER_0_110_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1__f__02687_ clknet_0__02687_ VGND VGND VPWR VPWR clknet_1_1__leaf__02687_
+ sky130_fd_sc_hd__clkbuf_16
X_14487__611 clknet_1_1__leaf__02665_ VGND VGND VPWR VPWR net643 sky130_fd_sc_hd__inv_2
XFILLER_0_86_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_08871_ _04571_ _04574_ VGND VGND VPWR VPWR _04591_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_4_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14227__402 clknet_1_1__leaf__08432_ VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__inv_2
XFILLER_0_126_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09423_ CPU.PC\[14\] _04923_ VGND VGND VPWR VPWR _05126_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09354_ _04252_ _04699_ _04808_ CPU.aluReg\[17\] _05059_ VGND VGND VPWR VPWR _05060_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_23_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09285_ _04343_ _04993_ VGND VGND VPWR VPWR _04994_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_134_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_151_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_15153__1180 clknet_1_0__leaf__02746_ VGND VGND VPWR VPWR net1212 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_54_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10060_ _05625_ VGND VGND VPWR VPWR _02387_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f__03963_ clknet_0__03963_ VGND VGND VPWR VPWR clknet_1_0__leaf__03963_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_98_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10962_ _06182_ VGND VGND VPWR VPWR _02027_ sky130_fd_sc_hd__clkbuf_1
X_13750_ _07274_ _08167_ VGND VGND VPWR VPWR _08168_ sky130_fd_sc_hd__or2_1
X_14700__804 clknet_1_0__leaf__02685_ VGND VGND VPWR VPWR net836 sky130_fd_sc_hd__inv_2
X_15254__161 clknet_1_1__leaf__02756_ VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__inv_2
X_12701_ net1423 _07182_ VGND VGND VPWR VPWR _07183_ sky130_fd_sc_hd__or2_1
X_13681_ CPU.registerFile\[5\]\[23\] _07373_ _08100_ _07368_ VGND VGND VPWR VPWR _08101_
+ sky130_fd_sc_hd__o211a_1
X_10893_ net1667 _05675_ _06143_ VGND VGND VPWR VPWR _06146_ sky130_fd_sc_hd__mux2_1
XFILLER_0_156_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15420_ _08397_ _02909_ _02913_ _02916_ VGND VGND VPWR VPWR _02917_ sky130_fd_sc_hd__o22a_1
X_12632_ CPU.cycles\[4\] _07138_ net1355 VGND VGND VPWR VPWR _07141_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_155_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_12563_ _07104_ VGND VGND VPWR VPWR _01277_ sky130_fd_sc_hd__clkbuf_1
X_15351_ _02760_ VGND VGND VPWR VPWR _02849_ sky130_fd_sc_hd__buf_4
XFILLER_0_65_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_136_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11514_ CPU.mem_rstrb _06468_ _04783_ net1336 VGND VGND VPWR VPWR _06479_ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18070_ net133 _02350_ VGND VGND VPWR VPWR CPU.registerFile\[18\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_12494_ net2227 _05706_ _07060_ VGND VGND VPWR VPWR _07068_ sky130_fd_sc_hd__mux2_1
X_15282_ CPU.registerFile\[9\]\[0\] _02778_ _02780_ VGND VGND VPWR VPWR _02781_ sky130_fd_sc_hd__o21a_1
X_17021_ net279 _01343_ VGND VGND VPWR VPWR CPU.registerFile\[3\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_11445_ _05501_ net2194 _06433_ VGND VGND VPWR VPWR _06439_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0__02710_ _02710_ VGND VGND VPWR VPWR clknet_0__02710_ sky130_fd_sc_hd__clkbuf_16
X_14164_ CPU.Bimm\[5\] _04776_ _08413_ VGND VGND VPWR VPWR _08419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_151_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_11376_ _06402_ VGND VGND VPWR VPWR _01833_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_156_Right_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_13115_ CPU.registerFile\[15\]\[6\] _07281_ _07521_ CPU.registerFile\[11\]\[6\] _07253_
+ VGND VGND VPWR VPWR _07552_ sky130_fd_sc_hd__o221a_1
X_10327_ _05784_ VGND VGND VPWR VPWR _02264_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14095_ _04716_ _05313_ _08374_ VGND VGND VPWR VPWR _08375_ sky130_fd_sc_hd__a21bo_1
X_13046_ _07418_ _07481_ _07484_ VGND VGND VPWR VPWR _07485_ sky130_fd_sc_hd__o21a_1
X_17923_ net1112 _02207_ VGND VGND VPWR VPWR mapped_spi_flash.cmd_addr\[3\] sky130_fd_sc_hd__dfxtp_1
X_10258_ _05747_ VGND VGND VPWR VPWR _02311_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17854_ net1043 _02138_ VGND VGND VPWR VPWR CPU.registerFile\[28\]\[12\] sky130_fd_sc_hd__dfxtp_1
X_10189_ _05089_ VGND VGND VPWR VPWR _05702_ sky130_fd_sc_hd__clkbuf_4
X_16805_ per_uart.uart0.txd_reg\[0\] _07179_ VGND VGND VPWR VPWR _04113_ sky130_fd_sc_hd__nor2_1
X_17785_ net974 _02069_ VGND VGND VPWR VPWR CPU.registerFile\[2\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_16736_ _03991_ net1972 VGND VGND VPWR VPWR _04056_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_85_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_13968__252 clknet_1_0__leaf__08357_ VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__inv_2
X_16667_ _03992_ _03997_ _06030_ VGND VGND VPWR VPWR _02582_ sky130_fd_sc_hd__a21oi_1
X_13879_ _07405_ _08289_ _08291_ _08292_ _07359_ VGND VGND VPWR VPWR _08293_ sky130_fd_sc_hd__a221o_1
XFILLER_0_158_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15618_ CPU.registerFile\[16\]\[6\] _02833_ _02836_ CPU.registerFile\[17\]\[6\] _02764_
+ VGND VGND VPWR VPWR _03111_ sky130_fd_sc_hd__o221a_1
XFILLER_0_9_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18337_ clknet_leaf_4_clk _02617_ VGND VGND VPWR VPWR per_uart.rx_data\[1\] sky130_fd_sc_hd__dfxtp_1
X_15549_ CPU.registerFile\[9\]\[5\] _02778_ _02780_ VGND VGND VPWR VPWR _03043_ sky130_fd_sc_hd__o21a_1
X_09070_ _04688_ VGND VGND VPWR VPWR _04783_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_142_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_18268_ clknet_leaf_1_clk _02548_ VGND VGND VPWR VPWR per_uart.uart0.rxd_reg\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_14222__398 clknet_1_0__leaf__08431_ VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__inv_2
XFILLER_0_71_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17219_ net409 _01507_ VGND VGND VPWR VPWR CPU.registerFile\[27\]\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18199_ net230 _02479_ VGND VGND VPWR VPWR CPU.registerFile\[15\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold702 CPU.registerFile\[28\]\[16\] VGND VGND VPWR VPWR net1943 sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 CPU.registerFile\[13\]\[24\] VGND VGND VPWR VPWR net1954 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold724 CPU.registerFile\[3\]\[0\] VGND VGND VPWR VPWR net1965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold735 CPU.registerFile\[15\]\[19\] VGND VGND VPWR VPWR net1976 sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 CPU.registerFile\[3\]\[26\] VGND VGND VPWR VPWR net1987 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold757 CPU.registerFile\[15\]\[14\] VGND VGND VPWR VPWR net1998 sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 CPU.registerFile\[24\]\[21\] VGND VGND VPWR VPWR net2009 sky130_fd_sc_hd__dlygate4sd3_1
X_09972_ _05578_ VGND VGND VPWR VPWR _02460_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_123_Right_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold779 CPU.registerFile\[16\]\[9\] VGND VGND VPWR VPWR net2020 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_08923_ _04642_ VGND VGND VPWR VPWR _04643_ sky130_fd_sc_hd__buf_6
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08854_ _04572_ _04573_ VGND VGND VPWR VPWR _04574_ sky130_fd_sc_hd__nand2_1
X_08785_ net2 VGND VGND VPWR VPWR _04505_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_28_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14541__660 clknet_1_0__leaf__02670_ VGND VGND VPWR VPWR net692 sky130_fd_sc_hd__inv_2
XFILLER_0_138_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_153_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09406_ net1939 _05109_ _04983_ VGND VGND VPWR VPWR _05110_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09337_ _04818_ _05042_ _05043_ _04916_ VGND VGND VPWR VPWR _05044_ sky130_fd_sc_hd__o22a_1
XFILLER_0_35_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_09268_ _04976_ _04977_ VGND VGND VPWR VPWR _04978_ sky130_fd_sc_hd__nand2_1
X_14459__587 clknet_1_1__leaf__02661_ VGND VGND VPWR VPWR net619 sky130_fd_sc_hd__inv_2
XFILLER_0_133_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09199_ CPU.Iimm\[3\] _04496_ _04820_ VGND VGND VPWR VPWR _04911_ sky130_fd_sc_hd__mux2_1
X_14197__375 clknet_1_0__leaf__08429_ VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__inv_2
XFILLER_0_43_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11230_ net1744 _05668_ _06324_ VGND VGND VPWR VPWR _06325_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_11161_ _06287_ VGND VGND VPWR VPWR _06288_ sky130_fd_sc_hd__buf_4
X_10112_ _05653_ VGND VGND VPWR VPWR _02363_ sky130_fd_sc_hd__clkbuf_1
X_11092_ _04662_ _06250_ VGND VGND VPWR VPWR _06251_ sky130_fd_sc_hd__nor2_2
X_10043_ _05616_ VGND VGND VPWR VPWR _02395_ sky130_fd_sc_hd__clkbuf_1
X_14851_ clknet_1_0__leaf__02697_ VGND VGND VPWR VPWR _02701_ sky130_fd_sc_hd__buf_1
Xhold73 mapped_spi_flash.div_counter\[1\] VGND VGND VPWR VPWR net1314 sky130_fd_sc_hd__dlygate4sd3_1
X_14624__735 clknet_1_1__leaf__02678_ VGND VGND VPWR VPWR net767 sky130_fd_sc_hd__inv_2
Xhold84 _02187_ VGND VGND VPWR VPWR net1325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 mapped_spi_ram.state\[2\] VGND VGND VPWR VPWR net1336 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ _08214_ _08217_ _07474_ VGND VGND VPWR VPWR _08218_ sky130_fd_sc_hd__a21oi_2
X_17570_ net759 _01858_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_11994_ _06765_ VGND VGND VPWR VPWR _01575_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_67_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_826 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_13733_ CPU.registerFile\[5\]\[25\] CPU.registerFile\[4\]\[25\] _07262_ VGND VGND
+ VPWR VPWR _08151_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10945_ net1793 _05727_ _06165_ VGND VGND VPWR VPWR _06173_ sky130_fd_sc_hd__mux2_1
X_16452_ CPU.registerFile\[21\]\[30\] CPU.registerFile\[23\]\[30\] _05440_ VGND VGND
+ VPWR VPWR _03921_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13664_ CPU.registerFile\[28\]\[23\] _07987_ VGND VGND VPWR VPWR _08084_ sky130_fd_sc_hd__or2_1
X_10876_ net1808 _05727_ _06128_ VGND VGND VPWR VPWR _06136_ sky130_fd_sc_hd__mux2_1
X_15403_ _02872_ VGND VGND VPWR VPWR _02901_ sky130_fd_sc_hd__clkbuf_4
X_12615_ _07131_ VGND VGND VPWR VPWR _00009_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_80_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16383_ CPU.registerFile\[22\]\[28\] CPU.registerFile\[23\]\[28\] _02829_ VGND VGND
+ VPWR VPWR _03854_ sky130_fd_sc_hd__mux2_1
X_13595_ net1890 _07229_ _08016_ _08017_ VGND VGND VPWR VPWR _01315_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_80_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18122_ net185 _02402_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[20\] sky130_fd_sc_hd__dfxtp_1
X_15334_ _02832_ VGND VGND VPWR VPWR _02833_ sky130_fd_sc_hd__clkbuf_4
X_12546_ _07095_ VGND VGND VPWR VPWR _01285_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_696 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_18053_ net1226 _02333_ VGND VGND VPWR VPWR CPU.registerFile\[1\]\[15\] sky130_fd_sc_hd__dfxtp_1
X_15265_ _05070_ VGND VGND VPWR VPWR _02764_ sky130_fd_sc_hd__buf_4
X_12477_ net1865 _05689_ _07049_ VGND VGND VPWR VPWR _07059_ sky130_fd_sc_hd__mux2_1
X_14670__777 clknet_1_1__leaf__02682_ VGND VGND VPWR VPWR net809 sky130_fd_sc_hd__inv_2
XANTENNA_4 _02763_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_17004_ clknet_leaf_11_clk net1499 VGND VGND VPWR VPWR CPU.state\[3\] sky130_fd_sc_hd__dfxtp_2
X_11428_ _06429_ VGND VGND VPWR VPWR _01808_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_14147_ CPU.Jimm\[18\] _08408_ _08387_ VGND VGND VPWR VPWR _08409_ sky130_fd_sc_hd__mux2_1
X_11359_ _06392_ VGND VGND VPWR VPWR _01840_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_17906_ net1095 _02190_ VGND VGND VPWR VPWR mapped_spi_flash.rcv_data\[24\] sky130_fd_sc_hd__dfxtp_1
X_13029_ CPU.registerFile\[21\]\[4\] _07362_ _07383_ CPU.registerFile\[17\]\[4\] _07467_
+ VGND VGND VPWR VPWR _07468_ sky130_fd_sc_hd__o221a_2
X_17837_ net1026 _02121_ VGND VGND VPWR VPWR CPU.registerFile\[30\]\[27\] sky130_fd_sc_hd__dfxtp_1
Xrebuffer16 net1258 VGND VGND VPWR VPWR net1257 sky130_fd_sc_hd__dlygate4sd1_1
X_08570_ CPU.aluIn1\[1\] VGND VGND VPWR VPWR _04290_ sky130_fd_sc_hd__inv_2
Xrebuffer27 net1269 VGND VGND VPWR VPWR net1268 sky130_fd_sc_hd__dlymetal6s2s_1
X_17768_ net957 _02052_ VGND VGND VPWR VPWR CPU.registerFile\[5\]\[22\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xrebuffer38 net1281 VGND VGND VPWR VPWR net1279 sky130_fd_sc_hd__clkbuf_2
X_14599__712 clknet_1_1__leaf__02676_ VGND VGND VPWR VPWR net744 sky130_fd_sc_hd__inv_2
Xrebuffer49 net1295 VGND VGND VPWR VPWR net1296 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_0_77_804 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16719_ _03995_ _05203_ _07132_ VGND VGND VPWR VPWR _04042_ sky130_fd_sc_hd__o21ai_1
X_17699_ net888 _01987_ VGND VGND VPWR VPWR CPU.registerFile\[7\]\[21\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_135_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09122_ CPU.PC\[19\] _04832_ VGND VGND VPWR VPWR _04834_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_09053_ _04354_ _04766_ _04374_ VGND VGND VPWR VPWR _04767_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_853 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_131_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold510 CPU.registerFile\[27\]\[14\] VGND VGND VPWR VPWR net1751 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold521 CPU.PC\[23\] VGND VGND VPWR VPWR net1762 sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 CPU.registerFile\[30\]\[8\] VGND VGND VPWR VPWR net1773 sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 CPU.registerFile\[14\]\[17\] VGND VGND VPWR VPWR net1784 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold554 CPU.registerFile\[24\]\[23\] VGND VGND VPWR VPWR net1795 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold565 CPU.registerFile\[31\]\[4\] VGND VGND VPWR VPWR net1806 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold576 CPU.registerFile\[16\]\[3\] VGND VGND VPWR VPWR net1817 sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 CPU.registerFile\[19\]\[26\] VGND VGND VPWR VPWR net1828 sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 per_uart.uart0.rx_bitcount\[2\] VGND VGND VPWR VPWR net1839 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_09955_ _05569_ VGND VGND VPWR VPWR _02468_ sky130_fd_sc_hd__clkbuf_1
X_08906_ _04528_ net1280 VGND VGND VPWR VPWR _04626_ sky130_fd_sc_hd__or2_1
X_09886_ _05525_ VGND VGND VPWR VPWR _02493_ sky130_fd_sc_hd__clkbuf_1
Xhold1210 CPU.registerFile\[15\]\[4\] VGND VGND VPWR VPWR net2451 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_146_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1221 CPU.registerFile\[21\]\[10\] VGND VGND VPWR VPWR net2462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1232 CPU.registerFile\[20\]\[26\] VGND VGND VPWR VPWR net2473 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1243 CPU.aluReg\[6\] VGND VGND VPWR VPWR net2484 sky130_fd_sc_hd__dlygate4sd3_1
X_08837_ CPU.aluIn1\[15\] CPU.aluIn1\[14\] _04494_ VGND VGND VPWR VPWR _04557_ sky130_fd_sc_hd__o21ai_1
Xhold1254 CPU.registerFile\[14\]\[6\] VGND VGND VPWR VPWR net2495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1265 CPU.registerFile\[7\]\[10\] VGND VGND VPWR VPWR net2506 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1276 CPU.aluReg\[4\] VGND VGND VPWR VPWR net2517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1287 CPU.registerFile\[4\]\[23\] VGND VGND VPWR VPWR net2528 sky130_fd_sc_hd__dlygate4sd3_1
X_08768_ _04483_ _04487_ VGND VGND VPWR VPWR _04488_ sky130_fd_sc_hd__and2_1
Xhold1298 net9 VGND VGND VPWR VPWR net2539 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_405 _03528_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_416 clknet_1_0__leaf__07219_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_08699_ _04308_ _04285_ VGND VGND VPWR VPWR _04419_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_656 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_10730_ _05537_ net2143 _06056_ VGND VGND VPWR VPWR _06059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_10661_ _06018_ VGND VGND VPWR VPWR _06019_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_62_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_12400_ _07018_ VGND VGND VPWR VPWR _01387_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13380_ CPU.registerFile\[1\]\[14\] _07387_ _07808_ _07379_ VGND VGND VPWR VPWR _07809_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_63_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_14205__382 clknet_1_0__leaf__08430_ VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__inv_2
X_14812__905 clknet_1_0__leaf__02696_ VGND VGND VPWR VPWR net937 sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_11_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10592_ net1475 _05968_ _05977_ _05936_ VGND VGND VPWR VPWR _02191_ sky130_fd_sc_hd__o211a_1
X_12331_ _04748_ net2228 _06977_ VGND VGND VPWR VPWR _06982_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_12752__205 clknet_1_1__leaf__07221_ VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__inv_2
X_12262_ CPU.aluReg\[14\] _06931_ _06924_ VGND VGND VPWR VPWR _06932_ sky130_fd_sc_hd__mux2_1
X_11213_ _06315_ VGND VGND VPWR VPWR _01909_ sky130_fd_sc_hd__clkbuf_1
Xoutput6 net6 VGND VGND VPWR VPWR TXD sky130_fd_sc_hd__clkbuf_4
X_12193_ CPU.aluReg\[30\] _06878_ _06862_ VGND VGND VPWR VPWR _06879_ sky130_fd_sc_hd__mux2_1
X_11144_ net2319 _05721_ _06274_ VGND VGND VPWR VPWR _06279_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_15952_ CPU.registerFile\[15\]\[16\] CPU.registerFile\[11\]\[16\] _02906_ VGND VGND
+ VPWR VPWR _03435_ sky130_fd_sc_hd__mux2_1
X_11075_ net2146 _05721_ _06237_ VGND VGND VPWR VPWR _06242_ sky130_fd_sc_hd__mux2_1
X_10026_ net2294 _04982_ _05607_ VGND VGND VPWR VPWR _05608_ sky130_fd_sc_hd__mux2_1
X_15883_ CPU.registerFile\[8\]\[14\] _02789_ _03117_ _03367_ VGND VGND VPWR VPWR _03368_
+ sky130_fd_sc_hd__o211a_1
X_17622_ net811 _01910_ VGND VGND VPWR VPWR CPU.registerFile\[22\]\[8\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_19_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_17553_ net742 _01841_ VGND VGND VPWR VPWR CPU.registerFile\[23\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11977_ _06756_ VGND VGND VPWR VPWR _01583_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_13716_ CPU.registerFile\[31\]\[24\] _07556_ _07557_ CPU.registerFile\[27\]\[24\]
+ _07345_ VGND VGND VPWR VPWR _08135_ sky130_fd_sc_hd__o221a_1
XFILLER_0_129_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_10928_ net1567 _05710_ _06154_ VGND VGND VPWR VPWR _06164_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_17484_ net673 _01772_ VGND VGND VPWR VPWR CPU.mem_wbusy sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_128_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_829 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_16435_ _02848_ _03899_ _03903_ _02903_ VGND VGND VPWR VPWR _03904_ sky130_fd_sc_hd__o211a_1
X_13647_ CPU.registerFile\[8\]\[22\] CPU.registerFile\[12\]\[22\] _07785_ VGND VGND
+ VPWR VPWR _08068_ sky130_fd_sc_hd__mux2_1
X_10859_ net2480 _05710_ _06117_ VGND VGND VPWR VPWR _06127_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16366_ _02797_ _03834_ _03835_ _03836_ _02807_ VGND VGND VPWR VPWR _03837_ sky130_fd_sc_hd__a221o_1
X_13578_ CPU.registerFile\[14\]\[20\] CPU.registerFile\[10\]\[20\] _07480_ VGND VGND
+ VPWR VPWR _08001_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_18105_ net168 _02385_ VGND VGND VPWR VPWR CPU.registerFile\[17\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_15317_ _08403_ VGND VGND VPWR VPWR _02816_ sky130_fd_sc_hd__buf_4
X_12529_ net1748 _04695_ _07085_ VGND VGND VPWR VPWR _07087_ sky130_fd_sc_hd__mux2_1
X_16297_ _03195_ _03767_ _03769_ _02965_ VGND VGND VPWR VPWR _03770_ sky130_fd_sc_hd__a211o_1
XFILLER_0_41_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_113_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_18036_ net1209 _02316_ VGND VGND VPWR VPWR CPU.registerFile\[20\]\[30\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_93_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_09740_ CPU.aluIn1\[0\] _04302_ _04698_ _04218_ CPU.aluReg\[0\] VGND VGND VPWR VPWR
+ _05429_ sky130_fd_sc_hd__a32o_1
X_14908__991 clknet_1_0__leaf__02706_ VGND VGND VPWR VPWR net1023 sky130_fd_sc_hd__inv_2

